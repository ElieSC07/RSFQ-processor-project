.subckt Control_Unit_final_route bit7t bit6t bit5t bit4t bit3t bit2t bit1t overflowt zerot negt GCLKt Imm3 Imm2 Imm1 Imm0 select1 select0 read Addr1 Addr0 write_flags Op_Arith Op_And Op_Xor Cmpl_b1 Cmpl_b0 Cin readNextInstr1 readNextInstr0 nextInstrAddr1_1 nextInstrAddr1_0 nextInstrAddr0_1 nextInstrAddr0_0

X696 X546-SPLITT-OUT-R-IN X546-SPLITT-OUT-R-INr LSmitll_PTLRX
X697 X546-SPLITT-OUT-R-INr X546-SPLITT-OUT-R-INdc LSmitll_SFQDC
R698 X546-SPLITT-OUT-R-INdc 0 5
X699 X546-SPLITT-OUT-R-IN PAD

X700 X547-SPLITT-OUT-R-IN X547-SPLITT-OUT-R-INr LSmitll_PTLRX
X701 X547-SPLITT-OUT-R-INr X547-SPLITT-OUT-R-INdc LSmitll_SFQDC
R702 X547-SPLITT-OUT-R-INdc 0 5
X703 X547-SPLITT-OUT-R-IN PAD

X704 X548-SPLITT-OUT-R-IN X548-SPLITT-OUT-R-INr LSmitll_PTLRX
X705 X548-SPLITT-OUT-R-INr X548-SPLITT-OUT-R-INdc LSmitll_SFQDC
R706 X548-SPLITT-OUT-R-INdc 0 5
X707 X548-SPLITT-OUT-R-IN PAD

X708 X549-SPLITT-OUT-R-IN X549-SPLITT-OUT-R-INr LSmitll_PTLRX
X709 X549-SPLITT-OUT-R-INr X549-SPLITT-OUT-R-INdc LSmitll_SFQDC
R710 X549-SPLITT-OUT-R-INdc 0 5
X711 X549-SPLITT-OUT-R-IN PAD

X712 X550-SPLITT-OUT-R-IN X550-SPLITT-OUT-R-INr LSmitll_PTLRX
X713 X550-SPLITT-OUT-R-INr X550-SPLITT-OUT-R-INdc LSmitll_SFQDC
R714 X550-SPLITT-OUT-R-INdc 0 5
X715 X550-SPLITT-OUT-R-IN PAD

X716 X551-SPLITT-OUT-R-IN X551-SPLITT-OUT-R-INr LSmitll_PTLRX
X717 X551-SPLITT-OUT-R-INr X551-SPLITT-OUT-R-INdc LSmitll_SFQDC
R718 X551-SPLITT-OUT-R-INdc 0 5
X719 X551-SPLITT-OUT-R-IN PAD

X720 X552-SPLITT-OUT-R-IN X552-SPLITT-OUT-R-INr LSmitll_PTLRX
X721 X552-SPLITT-OUT-R-INr X552-SPLITT-OUT-R-INdc LSmitll_SFQDC
R722 X552-SPLITT-OUT-R-INdc 0 5
X723 X552-SPLITT-OUT-R-IN PAD

X724 X553-SPLITT-OUT-R-IN X553-SPLITT-OUT-R-INr LSmitll_PTLRX
X725 X553-SPLITT-OUT-R-INr X553-SPLITT-OUT-R-INdc LSmitll_SFQDC
R726 X553-SPLITT-OUT-R-INdc 0 5
X727 X553-SPLITT-OUT-R-IN PAD

X728 X554-SPLITT-OUT-R-IN X554-SPLITT-OUT-R-INr LSmitll_PTLRX
X729 X554-SPLITT-OUT-R-INr X554-SPLITT-OUT-R-INdc LSmitll_SFQDC
R730 X554-SPLITT-OUT-R-INdc 0 5
X731 X554-SPLITT-OUT-R-IN PAD

X732 X555-SPLITT-OUT-R-IN X555-SPLITT-OUT-R-INr LSmitll_PTLRX
X733 X555-SPLITT-OUT-R-INr X555-SPLITT-OUT-R-INdc LSmitll_SFQDC
R734 X555-SPLITT-OUT-R-INdc 0 5
X735 X555-SPLITT-OUT-R-IN PAD

X736 X556-SPLITT-OUT-R-IN X556-SPLITT-OUT-R-INr LSmitll_PTLRX
X737 X556-SPLITT-OUT-R-INr X556-SPLITT-OUT-R-INdc LSmitll_SFQDC
R738 X556-SPLITT-OUT-R-INdc 0 5
X739 X556-SPLITT-OUT-R-IN PAD

X740 X557-SPLITT-OUT-R-IN X557-SPLITT-OUT-R-INr LSmitll_PTLRX
X741 X557-SPLITT-OUT-R-INr X557-SPLITT-OUT-R-INdc LSmitll_SFQDC
R742 X557-SPLITT-OUT-R-INdc 0 5
X743 X557-SPLITT-OUT-R-IN PAD

X744 X558-SPLITT-OUT-R-IN X558-SPLITT-OUT-R-INr LSmitll_PTLRX
X745 X558-SPLITT-OUT-R-INr X558-SPLITT-OUT-R-INdc LSmitll_SFQDC
R746 X558-SPLITT-OUT-R-INdc 0 5
X747 X558-SPLITT-OUT-R-IN PAD

X748 X559-SPLITT-OUT-R-IN X559-SPLITT-OUT-R-INr LSmitll_PTLRX
X749 X559-SPLITT-OUT-R-INr X559-SPLITT-OUT-R-INdc LSmitll_SFQDC
R750 X559-SPLITT-OUT-R-INdc 0 5
X751 X559-SPLITT-OUT-R-IN PAD

X752 X560-SPLITT-OUT-R-IN X560-SPLITT-OUT-R-INr LSmitll_PTLRX
X753 X560-SPLITT-OUT-R-INr X560-SPLITT-OUT-R-INdc LSmitll_SFQDC
R754 X560-SPLITT-OUT-R-INdc 0 5
X755 X560-SPLITT-OUT-R-IN PAD

X756 X561-SPLITT-OUT-R-IN X561-SPLITT-OUT-R-INr LSmitll_PTLRX
X757 X561-SPLITT-OUT-R-INr X561-SPLITT-OUT-R-INdc LSmitll_SFQDC
R758 X561-SPLITT-OUT-R-INdc 0 5
X759 X561-SPLITT-OUT-R-IN PAD

X760 X562-SPLITT-OUT-R-IN X562-SPLITT-OUT-R-INr LSmitll_PTLRX
X761 X562-SPLITT-OUT-R-INr X562-SPLITT-OUT-R-INdc LSmitll_SFQDC
R762 X562-SPLITT-OUT-R-INdc 0 5
X763 X562-SPLITT-OUT-R-IN PAD

X764 X563-SPLITT-OUT-R-IN X563-SPLITT-OUT-R-INr LSmitll_PTLRX
X765 X563-SPLITT-OUT-R-INr X563-SPLITT-OUT-R-INdc LSmitll_SFQDC
R766 X563-SPLITT-OUT-R-INdc 0 5
X767 X563-SPLITT-OUT-R-IN PAD

X768 X564-SPLITT-OUT-R-IN X564-SPLITT-OUT-R-INr LSmitll_PTLRX
X769 X564-SPLITT-OUT-R-INr X564-SPLITT-OUT-R-INdc LSmitll_SFQDC
R770 X564-SPLITT-OUT-R-INdc 0 5
X771 X564-SPLITT-OUT-R-IN PAD

X772 X565-SPLITT-OUT-R-IN X565-SPLITT-OUT-R-INr LSmitll_PTLRX
X773 X565-SPLITT-OUT-R-INr X565-SPLITT-OUT-R-INdc LSmitll_SFQDC
R774 X565-SPLITT-OUT-R-INdc 0 5
X775 X565-SPLITT-OUT-R-IN PAD

X776 X566-SPLITT-OUT-R-IN X566-SPLITT-OUT-R-INr LSmitll_PTLRX
X777 X566-SPLITT-OUT-R-INr X566-SPLITT-OUT-R-INdc LSmitll_SFQDC
R778 X566-SPLITT-OUT-R-INdc 0 5
X779 X566-SPLITT-OUT-R-IN PAD



t784 X1-LSmitll_SPLITT-OUT-X4-LSmitll_NOTT-INt 0 X1-LSmitll_SPLITT-OUT-X4-LSmitll_NOTT-IN 0 z0=5 td=3.5ps
t785 X1-LSmitll_SPLITT-OUT-X3-LSmitll_DFFT-INt 0 X1-LSmitll_SPLITT-OUT-X3-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X1 bit7 X1-LSmitll_SPLITT-OUT-X4-LSmitll_NOTT-INt X1-LSmitll_SPLITT-OUT-X3-LSmitll_DFFT-INt LSmitll_SPLITT

t786 X2-LSmitll_SPLITT-OUT-X6-LSmitll_NOTT-INt 0 X2-LSmitll_SPLITT-OUT-X6-LSmitll_NOTT-IN 0 z0=5 td=4.6ps
t787 X2-LSmitll_SPLITT-OUT-X5-LSmitll_DFFT-INt 0 X2-LSmitll_SPLITT-OUT-X5-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X2 bit6 X2-LSmitll_SPLITT-OUT-X6-LSmitll_NOTT-INt X2-LSmitll_SPLITT-OUT-X5-LSmitll_DFFT-INt LSmitll_SPLITT

t788 X3-LSmitll_DFFT-OUT-X21-LSmitll_SPLITT-INt 0 X3-LSmitll_DFFT-OUT-X21-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X3 X1-LSmitll_SPLITT-OUT-X3-LSmitll_DFFT-IN X452-LSmitll_SPLITT-OUT-X3-LSmitll_DFFT-IN X3-LSmitll_DFFT-OUT-X21-LSmitll_SPLITT-INt LSmitll_DFFT

t789 X4-LSmitll_NOTT-OUT-X20-LSmitll_SPLITT-INt 0 X4-LSmitll_NOTT-OUT-X20-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X4 X1-LSmitll_SPLITT-OUT-X4-LSmitll_NOTT-IN X546-LSmitll_SPLITT-OUT-X4-LSmitll_NOTT-IN X4-LSmitll_NOTT-OUT-X20-LSmitll_SPLITT-INt LSmitll_NOTT

t790 X5-LSmitll_DFFT-OUT-X23-LSmitll_SPLITT-INt 0 X5-LSmitll_DFFT-OUT-X23-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
X5 X2-LSmitll_SPLITT-OUT-X5-LSmitll_DFFT-IN X474-LSmitll_SPLITT-OUT-X5-LSmitll_DFFT-IN X5-LSmitll_DFFT-OUT-X23-LSmitll_SPLITT-INt LSmitll_DFFT

t791 X6-LSmitll_NOTT-OUT-X22-LSmitll_SPLITT-INt 0 X6-LSmitll_NOTT-OUT-X22-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X6 X2-LSmitll_SPLITT-OUT-X6-LSmitll_NOTT-IN X482-LSmitll_SPLITT-OUT-X6-LSmitll_NOTT-IN X6-LSmitll_NOTT-OUT-X22-LSmitll_SPLITT-INt LSmitll_NOTT

t792 X7-LSmitll_DFFT-OUT-X28-LSmitll_DFFT-INt 0 X7-LSmitll_DFFT-OUT-X28-LSmitll_DFFT-IN 0 z0=5 td=12.1ps
X7 bit5 X437-LSmitll_SPLITT-OUT-X7-LSmitll_DFFT-IN X7-LSmitll_DFFT-OUT-X28-LSmitll_DFFT-INt LSmitll_DFFT

t793 X8-LSmitll_DFFT-OUT-X29-LSmitll_DFFT-INt 0 X8-LSmitll_DFFT-OUT-X29-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X8 bit4 X434-LSmitll_SPLITT-OUT-X8-LSmitll_DFFT-IN X8-LSmitll_DFFT-OUT-X29-LSmitll_DFFT-INt LSmitll_DFFT

t794 X9-LSmitll_DFFT-OUT-X30-LSmitll_DFFT-INt 0 X9-LSmitll_DFFT-OUT-X30-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X9 bit3 X433-LSmitll_SPLITT-OUT-X9-LSmitll_DFFT-IN X9-LSmitll_DFFT-OUT-X30-LSmitll_DFFT-INt LSmitll_DFFT

t795 X10-LSmitll_DFFT-OUT-X31-LSmitll_DFFT-INt 0 X10-LSmitll_DFFT-OUT-X31-LSmitll_DFFT-IN 0 z0=5 td=4.0ps
X10 bit2 X459-LSmitll_SPLITT-OUT-X10-LSmitll_DFFT-IN X10-LSmitll_DFFT-OUT-X31-LSmitll_DFFT-INt LSmitll_DFFT

t796 X11-LSmitll_DFFT-OUT-X32-LSmitll_DFFT-INt 0 X11-LSmitll_DFFT-OUT-X32-LSmitll_DFFT-IN 0 z0=5 td=2.8ps
X11 bit1 X467-LSmitll_SPLITT-OUT-X11-LSmitll_DFFT-IN X11-LSmitll_DFFT-OUT-X32-LSmitll_DFFT-INt LSmitll_DFFT

t797 X12-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-INt 0 X12-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-IN 0 z0=5 td=2.3ps
t798 X12-LSmitll_SPLITT-OUT-X15-LSmitll_DFFT-INt 0 X12-LSmitll_SPLITT-OUT-X15-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X12 overflow X12-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-INt X12-LSmitll_SPLITT-OUT-X15-LSmitll_DFFT-INt LSmitll_SPLITT

t799 X13-LSmitll_SPLITT-OUT-X17-LSmitll_NOTT-INt 0 X13-LSmitll_SPLITT-OUT-X17-LSmitll_NOTT-IN 0 z0=5 td=3.3ps
t800 X13-LSmitll_SPLITT-OUT-X16-LSmitll_DFFT-INt 0 X13-LSmitll_SPLITT-OUT-X16-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X13 zero X13-LSmitll_SPLITT-OUT-X17-LSmitll_NOTT-INt X13-LSmitll_SPLITT-OUT-X16-LSmitll_DFFT-INt LSmitll_SPLITT

t801 X14-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-INt 0 X14-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-IN 0 z0=5 td=4.0ps
t802 X14-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-INt 0 X14-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X14 neg X14-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-INt X14-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-INt LSmitll_SPLITT

t803 X15-LSmitll_DFFT-OUT-X35-LSmitll_XORT-INt 0 X15-LSmitll_DFFT-OUT-X35-LSmitll_XORT-IN 0 z0=5 td=1.3ps
X15 X12-LSmitll_SPLITT-OUT-X15-LSmitll_DFFT-IN X430-LSmitll_SPLITT-OUT-X15-LSmitll_DFFT-IN X15-LSmitll_DFFT-OUT-X35-LSmitll_XORT-INt LSmitll_DFFT

t804 X16-LSmitll_DFFT-OUT-X33-LSmitll_DFFT-INt 0 X16-LSmitll_DFFT-OUT-X33-LSmitll_DFFT-IN 0 z0=5 td=26.7ps
X16 X13-LSmitll_SPLITT-OUT-X16-LSmitll_DFFT-IN X438-LSmitll_SPLITT-OUT-X16-LSmitll_DFFT-IN X16-LSmitll_DFFT-OUT-X33-LSmitll_DFFT-INt LSmitll_DFFT

t805 X17-LSmitll_NOTT-OUT-X34-LSmitll_DFFT-INt 0 X17-LSmitll_NOTT-OUT-X34-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X17 X13-LSmitll_SPLITT-OUT-X17-LSmitll_NOTT-IN X460-LSmitll_SPLITT-OUT-X17-LSmitll_NOTT-IN X17-LSmitll_NOTT-OUT-X34-LSmitll_DFFT-INt LSmitll_NOTT

t806 X18-LSmitll_DFFT-OUT-X35-LSmitll_XORT-INt 0 X18-LSmitll_DFFT-OUT-X35-LSmitll_XORT-IN 0 z0=5 td=2.3ps
X18 X14-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-IN X349-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-IN X18-LSmitll_DFFT-OUT-X35-LSmitll_XORT-INt LSmitll_DFFT

t807 X19-LSmitll_XORT-OUT-X36-LSmitll_NOTT-INt 0 X19-LSmitll_XORT-OUT-X36-LSmitll_NOTT-IN 0 z0=5 td=3.9ps
X19 X12-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-IN X14-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-IN X431-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-IN X19-LSmitll_XORT-OUT-X36-LSmitll_NOTT-INt LSmitll_XORT

t808 X20-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-INt 0 X20-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-IN 0 z0=5 td=4.3ps
t809 X20-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-INt 0 X20-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X20 X4-LSmitll_NOTT-OUT-X20-LSmitll_SPLITT-IN X20-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-INt X20-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-INt LSmitll_SPLITT

t810 X21-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-INt 0 X21-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
t811 X21-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-INt 0 X21-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-IN 0 z0=5 td=3.9ps
X21 X3-LSmitll_DFFT-OUT-X21-LSmitll_SPLITT-IN X21-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-INt X21-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-INt LSmitll_SPLITT

t812 X22-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-INt 0 X22-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-IN 0 z0=5 td=5.4ps
t813 X22-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-INt 0 X22-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
X22 X6-LSmitll_NOTT-OUT-X22-LSmitll_SPLITT-IN X22-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-INt X22-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-INt LSmitll_SPLITT

t814 X23-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-INt 0 X23-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-IN 0 z0=5 td=3.9ps
t815 X23-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-INt 0 X23-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
X23 X5-LSmitll_DFFT-OUT-X23-LSmitll_SPLITT-IN X23-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-INt X23-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-INt LSmitll_SPLITT

t816 X24-LSmitll_AND2T-OUT-X68-LSmitll_DFFT-INt 0 X24-LSmitll_AND2T-OUT-X68-LSmitll_DFFT-IN 0 z0=5 td=29.5ps
X24 X20-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-IN X22-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-IN X482-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-IN X24-LSmitll_AND2T-OUT-X68-LSmitll_DFFT-INt LSmitll_AND2T

t817 X25-LSmitll_AND2T-OUT-X43-LSmitll_SPLITT-INt 0 X25-LSmitll_AND2T-OUT-X43-LSmitll_SPLITT-IN 0 z0=5 td=20.3ps
X25 X20-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-IN X23-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-IN X547-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-IN X25-LSmitll_AND2T-OUT-X43-LSmitll_SPLITT-INt LSmitll_AND2T

t818 X26-LSmitll_AND2T-OUT-X44-LSmitll_SPLITT-INt 0 X26-LSmitll_AND2T-OUT-X44-LSmitll_SPLITT-IN 0 z0=5 td=4.3ps
X26 X22-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-IN X21-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-IN X476-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-IN X26-LSmitll_AND2T-OUT-X44-LSmitll_SPLITT-INt LSmitll_AND2T

t819 X27-LSmitll_AND2T-OUT-X40-LSmitll_SPLITT-INt 0 X27-LSmitll_AND2T-OUT-X40-LSmitll_SPLITT-IN 0 z0=5 td=11.6ps
X27 X21-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-IN X23-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-IN X454-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-IN X27-LSmitll_AND2T-OUT-X40-LSmitll_SPLITT-INt LSmitll_AND2T

t820 X28-LSmitll_DFFT-OUT-X45-LSmitll_SPLITT-INt 0 X28-LSmitll_DFFT-OUT-X45-LSmitll_SPLITT-IN 0 z0=5 td=8.4ps
X28 X7-LSmitll_DFFT-OUT-X28-LSmitll_DFFT-IN X345-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-IN X28-LSmitll_DFFT-OUT-X45-LSmitll_SPLITT-INt LSmitll_DFFT

t821 X29-LSmitll_DFFT-OUT-X48-LSmitll_SPLITT-INt 0 X29-LSmitll_DFFT-OUT-X48-LSmitll_SPLITT-IN 0 z0=5 td=12.3ps
X29 X8-LSmitll_DFFT-OUT-X29-LSmitll_DFFT-IN X433-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-IN X29-LSmitll_DFFT-OUT-X48-LSmitll_SPLITT-INt LSmitll_DFFT

t822 X30-LSmitll_DFFT-OUT-X51-LSmitll_SPLITT-INt 0 X30-LSmitll_DFFT-OUT-X51-LSmitll_SPLITT-IN 0 z0=5 td=6.1ps
X30 X9-LSmitll_DFFT-OUT-X30-LSmitll_DFFT-IN X548-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-IN X30-LSmitll_DFFT-OUT-X51-LSmitll_SPLITT-INt LSmitll_DFFT

t823 X31-LSmitll_DFFT-OUT-X52-LSmitll_SPLITT-INt 0 X31-LSmitll_DFFT-OUT-X52-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X31 X10-LSmitll_DFFT-OUT-X31-LSmitll_DFFT-IN X438-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-IN X31-LSmitll_DFFT-OUT-X52-LSmitll_SPLITT-INt LSmitll_DFFT

t824 X32-LSmitll_DFFT-OUT-X57-LSmitll_SPLITT-INt 0 X32-LSmitll_DFFT-OUT-X57-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X32 X11-LSmitll_DFFT-OUT-X32-LSmitll_DFFT-IN X467-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-IN X32-LSmitll_DFFT-OUT-X57-LSmitll_SPLITT-INt LSmitll_DFFT

t825 X33-LSmitll_DFFT-OUT-X37-LSmitll_SPLITT-INt 0 X33-LSmitll_DFFT-OUT-X37-LSmitll_SPLITT-IN 0 z0=5 td=5.4ps
X33 X16-LSmitll_DFFT-OUT-X33-LSmitll_DFFT-IN X320-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-IN X33-LSmitll_DFFT-OUT-X37-LSmitll_SPLITT-INt LSmitll_DFFT

t826 X34-LSmitll_DFFT-OUT-X90-LSmitll_AND2T-INt 0 X34-LSmitll_DFFT-OUT-X90-LSmitll_AND2T-IN 0 z0=5 td=22.3ps
X34 X17-LSmitll_NOTT-OUT-X34-LSmitll_DFFT-IN X466-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-IN X34-LSmitll_DFFT-OUT-X90-LSmitll_AND2T-INt LSmitll_DFFT

t827 X35-LSmitll_XORT-OUT-X39-LSmitll_SPLITT-INt 0 X35-LSmitll_XORT-OUT-X39-LSmitll_SPLITT-IN 0 z0=5 td=20.5ps
X35 X15-LSmitll_DFFT-OUT-X35-LSmitll_XORT-IN X18-LSmitll_DFFT-OUT-X35-LSmitll_XORT-IN X350-LSmitll_SPLITT-OUT-X35-LSmitll_XORT-IN X35-LSmitll_XORT-OUT-X39-LSmitll_SPLITT-INt LSmitll_XORT

t828 X36-LSmitll_NOTT-OUT-X38-LSmitll_SPLITT-INt 0 X36-LSmitll_NOTT-OUT-X38-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X36 X19-LSmitll_XORT-OUT-X36-LSmitll_NOTT-IN X437-LSmitll_SPLITT-OUT-X36-LSmitll_NOTT-IN X36-LSmitll_NOTT-OUT-X38-LSmitll_SPLITT-INt LSmitll_NOTT

t829 X37-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-INt 0 X37-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-IN 0 z0=5 td=1.7ps
t830 X37-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-INt 0 X37-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
X37 X33-LSmitll_DFFT-OUT-X37-LSmitll_SPLITT-IN X37-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-INt X37-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-INt LSmitll_SPLITT

t831 X38-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-INt 0 X38-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-IN 0 z0=5 td=2.5ps
t832 X38-LSmitll_SPLITT-OUT-X90-LSmitll_AND2T-INt 0 X38-LSmitll_SPLITT-OUT-X90-LSmitll_AND2T-IN 0 z0=5 td=3.5ps
X38 X36-LSmitll_NOTT-OUT-X38-LSmitll_SPLITT-IN X38-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-INt X38-LSmitll_SPLITT-OUT-X90-LSmitll_AND2T-INt LSmitll_SPLITT

t833 X39-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-INt 0 X39-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-IN 0 z0=5 td=1.8ps
t834 X39-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-INt 0 X39-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X39 X35-LSmitll_XORT-OUT-X39-LSmitll_SPLITT-IN X39-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-INt X39-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-INt LSmitll_SPLITT

t835 X40-LSmitll_SPLITT-OUT-X42-LSmitll_SPLITT-INt 0 X40-LSmitll_SPLITT-OUT-X42-LSmitll_SPLITT-IN 0 z0=5 td=4.3ps
t836 X40-LSmitll_SPLITT-OUT-X41-LSmitll_SPLITT-INt 0 X40-LSmitll_SPLITT-OUT-X41-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X40 X27-LSmitll_AND2T-OUT-X40-LSmitll_SPLITT-IN X40-LSmitll_SPLITT-OUT-X42-LSmitll_SPLITT-INt X40-LSmitll_SPLITT-OUT-X41-LSmitll_SPLITT-INt LSmitll_SPLITT

t837 X41-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-INt 0 X41-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t838 X41-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-INt 0 X41-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
X41 X40-LSmitll_SPLITT-OUT-X41-LSmitll_SPLITT-IN X41-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-INt X41-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-INt LSmitll_SPLITT

t839 X42-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-INt 0 X42-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
t840 X42-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-INt 0 X42-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-IN 0 z0=5 td=5.6ps
X42 X40-LSmitll_SPLITT-OUT-X42-LSmitll_SPLITT-IN X42-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-INt X42-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-INt LSmitll_SPLITT

t841 X43-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-INt 0 X43-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
t842 X43-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-INt 0 X43-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-IN 0 z0=5 td=4.8ps
X43 X25-LSmitll_AND2T-OUT-X43-LSmitll_SPLITT-IN X43-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-INt X43-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-INt LSmitll_SPLITT

t843 X44-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-INt 0 X44-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-IN 0 z0=5 td=5.1ps
t844 X44-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-INt 0 X44-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-IN 0 z0=5 td=4.0ps
X44 X26-LSmitll_AND2T-OUT-X44-LSmitll_SPLITT-IN X44-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-INt X44-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-INt LSmitll_SPLITT

t845 X45-LSmitll_SPLITT-OUT-X47-LSmitll_SPLITT-INt 0 X45-LSmitll_SPLITT-OUT-X47-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t846 X45-LSmitll_SPLITT-OUT-X46-LSmitll_SPLITT-INt 0 X45-LSmitll_SPLITT-OUT-X46-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X45 X28-LSmitll_DFFT-OUT-X45-LSmitll_SPLITT-IN X45-LSmitll_SPLITT-OUT-X47-LSmitll_SPLITT-INt X45-LSmitll_SPLITT-OUT-X46-LSmitll_SPLITT-INt LSmitll_SPLITT

t847 X46-LSmitll_SPLITT-OUT-X70-LSmitll_DFFT-INt 0 X46-LSmitll_SPLITT-OUT-X70-LSmitll_DFFT-IN 0 z0=5 td=6.0ps
t848 X46-LSmitll_SPLITT-OUT-X69-LSmitll_NOTT-INt 0 X46-LSmitll_SPLITT-OUT-X69-LSmitll_NOTT-IN 0 z0=5 td=2.1ps
X46 X45-LSmitll_SPLITT-OUT-X46-LSmitll_SPLITT-IN X46-LSmitll_SPLITT-OUT-X70-LSmitll_DFFT-INt X46-LSmitll_SPLITT-OUT-X69-LSmitll_NOTT-INt LSmitll_SPLITT

t849 X47-LSmitll_SPLITT-OUT-X72-LSmitll_DFFT-INt 0 X47-LSmitll_SPLITT-OUT-X72-LSmitll_DFFT-IN 0 z0=5 td=3.9ps
t850 X47-LSmitll_SPLITT-OUT-X71-LSmitll_DFFT-INt 0 X47-LSmitll_SPLITT-OUT-X71-LSmitll_DFFT-IN 0 z0=5 td=6.4ps
X47 X45-LSmitll_SPLITT-OUT-X47-LSmitll_SPLITT-IN X47-LSmitll_SPLITT-OUT-X72-LSmitll_DFFT-INt X47-LSmitll_SPLITT-OUT-X71-LSmitll_DFFT-INt LSmitll_SPLITT

t851 X48-LSmitll_SPLITT-OUT-X50-LSmitll_SPLITT-INt 0 X48-LSmitll_SPLITT-OUT-X50-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t852 X48-LSmitll_SPLITT-OUT-X49-LSmitll_SPLITT-INt 0 X48-LSmitll_SPLITT-OUT-X49-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X48 X29-LSmitll_DFFT-OUT-X48-LSmitll_SPLITT-IN X48-LSmitll_SPLITT-OUT-X50-LSmitll_SPLITT-INt X48-LSmitll_SPLITT-OUT-X49-LSmitll_SPLITT-INt LSmitll_SPLITT

t853 X49-LSmitll_SPLITT-OUT-X74-LSmitll_DFFT-INt 0 X49-LSmitll_SPLITT-OUT-X74-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
t854 X49-LSmitll_SPLITT-OUT-X73-LSmitll_DFFT-INt 0 X49-LSmitll_SPLITT-OUT-X73-LSmitll_DFFT-IN 0 z0=5 td=7.0ps
X49 X48-LSmitll_SPLITT-OUT-X49-LSmitll_SPLITT-IN X49-LSmitll_SPLITT-OUT-X74-LSmitll_DFFT-INt X49-LSmitll_SPLITT-OUT-X73-LSmitll_DFFT-INt LSmitll_SPLITT

t855 X50-LSmitll_SPLITT-OUT-X76-LSmitll_DFFT-INt 0 X50-LSmitll_SPLITT-OUT-X76-LSmitll_DFFT-IN 0 z0=5 td=4.4ps
t856 X50-LSmitll_SPLITT-OUT-X75-LSmitll_DFFT-INt 0 X50-LSmitll_SPLITT-OUT-X75-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X50 X48-LSmitll_SPLITT-OUT-X50-LSmitll_SPLITT-IN X50-LSmitll_SPLITT-OUT-X76-LSmitll_DFFT-INt X50-LSmitll_SPLITT-OUT-X75-LSmitll_DFFT-INt LSmitll_SPLITT

t857 X51-LSmitll_SPLITT-OUT-X55-LSmitll_SPLITT-INt 0 X51-LSmitll_SPLITT-OUT-X55-LSmitll_SPLITT-IN 0 z0=5 td=3.2ps
t858 X51-LSmitll_SPLITT-OUT-X53-LSmitll_SPLITT-INt 0 X51-LSmitll_SPLITT-OUT-X53-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
X51 X30-LSmitll_DFFT-OUT-X51-LSmitll_SPLITT-IN X51-LSmitll_SPLITT-OUT-X55-LSmitll_SPLITT-INt X51-LSmitll_SPLITT-OUT-X53-LSmitll_SPLITT-INt LSmitll_SPLITT

t859 X52-LSmitll_SPLITT-OUT-X56-LSmitll_SPLITT-INt 0 X52-LSmitll_SPLITT-OUT-X56-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t860 X52-LSmitll_SPLITT-OUT-X54-LSmitll_SPLITT-INt 0 X52-LSmitll_SPLITT-OUT-X54-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X52 X31-LSmitll_DFFT-OUT-X52-LSmitll_SPLITT-IN X52-LSmitll_SPLITT-OUT-X56-LSmitll_SPLITT-INt X52-LSmitll_SPLITT-OUT-X54-LSmitll_SPLITT-INt LSmitll_SPLITT

t861 X53-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-INt 0 X53-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
t862 X53-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-INt 0 X53-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X53 X51-LSmitll_SPLITT-OUT-X53-LSmitll_SPLITT-IN X53-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-INt X53-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-INt LSmitll_SPLITT

t863 X54-LSmitll_SPLITT-OUT-X82-LSmitll_DFFT-INt 0 X54-LSmitll_SPLITT-OUT-X82-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
t864 X54-LSmitll_SPLITT-OUT-X81-LSmitll_DFFT-INt 0 X54-LSmitll_SPLITT-OUT-X81-LSmitll_DFFT-IN 0 z0=5 td=4.7ps
X54 X52-LSmitll_SPLITT-OUT-X54-LSmitll_SPLITT-IN X54-LSmitll_SPLITT-OUT-X82-LSmitll_DFFT-INt X54-LSmitll_SPLITT-OUT-X81-LSmitll_DFFT-INt LSmitll_SPLITT

t865 X55-LSmitll_SPLITT-OUT-X80-LSmitll_NOTT-INt 0 X55-LSmitll_SPLITT-OUT-X80-LSmitll_NOTT-IN 0 z0=5 td=4.2ps
t866 X55-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-INt 0 X55-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X55 X51-LSmitll_SPLITT-OUT-X55-LSmitll_SPLITT-IN X55-LSmitll_SPLITT-OUT-X80-LSmitll_NOTT-INt X55-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-INt LSmitll_SPLITT

t867 X56-LSmitll_SPLITT-OUT-X84-LSmitll_NOTT-INt 0 X56-LSmitll_SPLITT-OUT-X84-LSmitll_NOTT-IN 0 z0=5 td=1.2ps
t868 X56-LSmitll_SPLITT-OUT-X83-LSmitll_DFFT-INt 0 X56-LSmitll_SPLITT-OUT-X83-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
X56 X52-LSmitll_SPLITT-OUT-X56-LSmitll_SPLITT-IN X56-LSmitll_SPLITT-OUT-X84-LSmitll_NOTT-INt X56-LSmitll_SPLITT-OUT-X83-LSmitll_DFFT-INt LSmitll_SPLITT

t869 X57-LSmitll_SPLITT-OUT-X59-LSmitll_SPLITT-INt 0 X57-LSmitll_SPLITT-OUT-X59-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t870 X57-LSmitll_SPLITT-OUT-X58-LSmitll_SPLITT-INt 0 X57-LSmitll_SPLITT-OUT-X58-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X57 X32-LSmitll_DFFT-OUT-X57-LSmitll_SPLITT-IN X57-LSmitll_SPLITT-OUT-X59-LSmitll_SPLITT-INt X57-LSmitll_SPLITT-OUT-X58-LSmitll_SPLITT-INt LSmitll_SPLITT

t871 X58-LSmitll_SPLITT-OUT-X86-LSmitll_DFFT-INt 0 X58-LSmitll_SPLITT-OUT-X86-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
t872 X58-LSmitll_SPLITT-OUT-X85-LSmitll_DFFT-INt 0 X58-LSmitll_SPLITT-OUT-X85-LSmitll_DFFT-IN 0 z0=5 td=4.2ps
X58 X57-LSmitll_SPLITT-OUT-X58-LSmitll_SPLITT-IN X58-LSmitll_SPLITT-OUT-X86-LSmitll_DFFT-INt X58-LSmitll_SPLITT-OUT-X85-LSmitll_DFFT-INt LSmitll_SPLITT

t873 X59-LSmitll_SPLITT-OUT-X88-LSmitll_NOTT-INt 0 X59-LSmitll_SPLITT-OUT-X88-LSmitll_NOTT-IN 0 z0=5 td=1.2ps
t874 X59-LSmitll_SPLITT-OUT-X87-LSmitll_DFFT-INt 0 X59-LSmitll_SPLITT-OUT-X87-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
X59 X57-LSmitll_SPLITT-OUT-X59-LSmitll_SPLITT-IN X59-LSmitll_SPLITT-OUT-X88-LSmitll_NOTT-INt X59-LSmitll_SPLITT-OUT-X87-LSmitll_DFFT-INt LSmitll_SPLITT

t875 X60-LSmitll_DFFT-OUT-X104-LSmitll_SPLITT-INt 0 X60-LSmitll_DFFT-OUT-X104-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X60 X41-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-IN X447-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-IN X60-LSmitll_DFFT-OUT-X104-LSmitll_SPLITT-INt LSmitll_DFFT

t876 X61-LSmitll_DFFT-OUT-X105-LSmitll_SPLITT-INt 0 X61-LSmitll_DFFT-OUT-X105-LSmitll_SPLITT-IN 0 z0=5 td=6.2ps
X61 X41-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-IN X448-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-IN X61-LSmitll_DFFT-OUT-X105-LSmitll_SPLITT-INt LSmitll_DFFT

t877 X62-LSmitll_DFFT-OUT-X106-LSmitll_SPLITT-INt 0 X62-LSmitll_DFFT-OUT-X106-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X62 X42-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-IN X359-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-IN X62-LSmitll_DFFT-OUT-X106-LSmitll_SPLITT-INt LSmitll_DFFT

t878 X63-LSmitll_DFFT-OUT-X107-LSmitll_SPLITT-INt 0 X63-LSmitll_DFFT-OUT-X107-LSmitll_SPLITT-IN 0 z0=5 td=9.9ps
X63 X42-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-IN X407-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-IN X63-LSmitll_DFFT-OUT-X107-LSmitll_SPLITT-INt LSmitll_DFFT

t879 X64-LSmitll_DFFT-OUT-X99-LSmitll_SPLITT-INt 0 X64-LSmitll_DFFT-OUT-X99-LSmitll_SPLITT-IN 0 z0=5 td=4.6ps
X64 X43-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-IN X401-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-IN X64-LSmitll_DFFT-OUT-X99-LSmitll_SPLITT-INt LSmitll_DFFT

t880 X65-LSmitll_DFFT-OUT-X102-LSmitll_SPLITT-INt 0 X65-LSmitll_DFFT-OUT-X102-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
X65 X43-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-IN X495-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-IN X65-LSmitll_DFFT-OUT-X102-LSmitll_SPLITT-INt LSmitll_DFFT

t881 X66-LSmitll_DFFT-OUT-X94-LSmitll_SPLITT-INt 0 X66-LSmitll_DFFT-OUT-X94-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
X66 X44-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-IN X451-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-IN X66-LSmitll_DFFT-OUT-X94-LSmitll_SPLITT-INt LSmitll_DFFT

t882 X67-LSmitll_DFFT-OUT-X97-LSmitll_SPLITT-INt 0 X67-LSmitll_DFFT-OUT-X97-LSmitll_SPLITT-IN 0 z0=5 td=10.3ps
X67 X44-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-IN X492-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-IN X67-LSmitll_DFFT-OUT-X97-LSmitll_SPLITT-INt LSmitll_DFFT

t883 X68-LSmitll_DFFT-OUT-X115-LSmitll_DFFT-INt 0 X68-LSmitll_DFFT-OUT-X115-LSmitll_DFFT-IN 0 z0=5 td=2.0ps
X68 X24-LSmitll_AND2T-OUT-X68-LSmitll_DFFT-IN X549-LSmitll_SPLITT-OUT-X68-LSmitll_DFFT-IN X68-LSmitll_DFFT-OUT-X115-LSmitll_DFFT-INt LSmitll_DFFT

t884 X69-LSmitll_NOTT-OUT-X109-LSmitll_SPLITT-INt 0 X69-LSmitll_NOTT-OUT-X109-LSmitll_SPLITT-IN 0 z0=5 td=4.4ps
X69 X46-LSmitll_SPLITT-OUT-X69-LSmitll_NOTT-IN X357-LSmitll_SPLITT-OUT-X69-LSmitll_NOTT-IN X69-LSmitll_NOTT-OUT-X109-LSmitll_SPLITT-INt LSmitll_NOTT

t885 X70-LSmitll_DFFT-OUT-X110-LSmitll_SPLITT-INt 0 X70-LSmitll_DFFT-OUT-X110-LSmitll_SPLITT-IN 0 z0=5 td=20.6ps
X70 X46-LSmitll_SPLITT-OUT-X70-LSmitll_DFFT-IN X362-LSmitll_SPLITT-OUT-X70-LSmitll_DFFT-IN X70-LSmitll_DFFT-OUT-X110-LSmitll_SPLITT-INt LSmitll_DFFT

t886 X71-LSmitll_DFFT-OUT-X135-LSmitll_OR2T-INt 0 X71-LSmitll_DFFT-OUT-X135-LSmitll_OR2T-IN 0 z0=5 td=0.9ps
X71 X47-LSmitll_SPLITT-OUT-X71-LSmitll_DFFT-IN X337-LSmitll_SPLITT-OUT-X71-LSmitll_DFFT-IN X71-LSmitll_DFFT-OUT-X135-LSmitll_OR2T-INt LSmitll_DFFT

t887 X72-LSmitll_DFFT-OUT-X142-LSmitll_DFFT-INt 0 X72-LSmitll_DFFT-OUT-X142-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X72 X47-LSmitll_SPLITT-OUT-X72-LSmitll_DFFT-IN X400-LSmitll_SPLITT-OUT-X72-LSmitll_DFFT-IN X72-LSmitll_DFFT-OUT-X142-LSmitll_DFFT-INt LSmitll_DFFT

t888 X73-LSmitll_DFFT-OUT-X125-LSmitll_AND2T-INt 0 X73-LSmitll_DFFT-OUT-X125-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
X73 X49-LSmitll_SPLITT-OUT-X73-LSmitll_DFFT-IN X334-LSmitll_SPLITT-OUT-X73-LSmitll_DFFT-IN X73-LSmitll_DFFT-OUT-X125-LSmitll_AND2T-INt LSmitll_DFFT

t889 X74-LSmitll_DFFT-OUT-X111-LSmitll_SPLITT-INt 0 X74-LSmitll_DFFT-OUT-X111-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X74 X49-LSmitll_SPLITT-OUT-X74-LSmitll_DFFT-IN X335-LSmitll_SPLITT-OUT-X74-LSmitll_DFFT-IN X74-LSmitll_DFFT-OUT-X111-LSmitll_SPLITT-INt LSmitll_DFFT

t890 X75-LSmitll_DFFT-OUT-X135-LSmitll_OR2T-INt 0 X75-LSmitll_DFFT-OUT-X135-LSmitll_OR2T-IN 0 z0=5 td=3.6ps
X75 X50-LSmitll_SPLITT-OUT-X75-LSmitll_DFFT-IN X330-LSmitll_SPLITT-OUT-X75-LSmitll_DFFT-IN X75-LSmitll_DFFT-OUT-X135-LSmitll_OR2T-INt LSmitll_DFFT

t891 X76-LSmitll_DFFT-OUT-X143-LSmitll_DFFT-INt 0 X76-LSmitll_DFFT-OUT-X143-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X76 X50-LSmitll_SPLITT-OUT-X76-LSmitll_DFFT-IN X379-LSmitll_SPLITT-OUT-X76-LSmitll_DFFT-IN X76-LSmitll_DFFT-OUT-X143-LSmitll_DFFT-INt LSmitll_DFFT

t892 X77-LSmitll_DFFT-OUT-X128-LSmitll_AND2T-INt 0 X77-LSmitll_DFFT-OUT-X128-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
X77 X53-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-IN X362-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-IN X77-LSmitll_DFFT-OUT-X128-LSmitll_AND2T-INt LSmitll_DFFT

t893 X78-LSmitll_DFFT-OUT-X112-LSmitll_SPLITT-INt 0 X78-LSmitll_DFFT-OUT-X112-LSmitll_SPLITT-IN 0 z0=5 td=6.9ps
X78 X53-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-IN X359-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-IN X78-LSmitll_DFFT-OUT-X112-LSmitll_SPLITT-INt LSmitll_DFFT

t894 X79-LSmitll_DFFT-OUT-X136-LSmitll_DFFT-INt 0 X79-LSmitll_DFFT-OUT-X136-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X79 X55-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-IN X320-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-IN X79-LSmitll_DFFT-OUT-X136-LSmitll_DFFT-INt LSmitll_DFFT

t895 X80-LSmitll_NOTT-OUT-X137-LSmitll_AND2T-INt 0 X80-LSmitll_NOTT-OUT-X137-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X80 X55-LSmitll_SPLITT-OUT-X80-LSmitll_NOTT-IN X316-LSmitll_SPLITT-OUT-X80-LSmitll_NOTT-IN X80-LSmitll_NOTT-OUT-X137-LSmitll_AND2T-INt LSmitll_NOTT

t896 X81-LSmitll_DFFT-OUT-X131-LSmitll_AND2T-INt 0 X81-LSmitll_DFFT-OUT-X131-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
X81 X54-LSmitll_SPLITT-OUT-X81-LSmitll_DFFT-IN X503-LSmitll_SPLITT-OUT-X81-LSmitll_DFFT-IN X81-LSmitll_DFFT-OUT-X131-LSmitll_AND2T-INt LSmitll_DFFT

t897 X82-LSmitll_DFFT-OUT-X113-LSmitll_SPLITT-INt 0 X82-LSmitll_DFFT-OUT-X113-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X82 X54-LSmitll_SPLITT-OUT-X82-LSmitll_DFFT-IN X550-LSmitll_SPLITT-OUT-X82-LSmitll_DFFT-IN X82-LSmitll_DFFT-OUT-X113-LSmitll_SPLITT-INt LSmitll_DFFT

t898 X83-LSmitll_DFFT-OUT-X138-LSmitll_AND2T-INt 0 X83-LSmitll_DFFT-OUT-X138-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X83 X56-LSmitll_SPLITT-OUT-X83-LSmitll_DFFT-IN X431-LSmitll_SPLITT-OUT-X83-LSmitll_DFFT-IN X83-LSmitll_DFFT-OUT-X138-LSmitll_AND2T-INt LSmitll_DFFT

t899 X84-LSmitll_NOTT-OUT-X139-LSmitll_AND2T-INt 0 X84-LSmitll_NOTT-OUT-X139-LSmitll_AND2T-IN 0 z0=5 td=16.9ps
X84 X56-LSmitll_SPLITT-OUT-X84-LSmitll_NOTT-IN X434-LSmitll_SPLITT-OUT-X84-LSmitll_NOTT-IN X84-LSmitll_NOTT-OUT-X139-LSmitll_AND2T-INt LSmitll_NOTT

t900 X85-LSmitll_DFFT-OUT-X134-LSmitll_AND2T-INt 0 X85-LSmitll_DFFT-OUT-X134-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
X85 X58-LSmitll_SPLITT-OUT-X85-LSmitll_DFFT-IN X530-LSmitll_SPLITT-OUT-X85-LSmitll_DFFT-IN X85-LSmitll_DFFT-OUT-X134-LSmitll_AND2T-INt LSmitll_DFFT

t901 X86-LSmitll_DFFT-OUT-X114-LSmitll_SPLITT-INt 0 X86-LSmitll_DFFT-OUT-X114-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X86 X58-LSmitll_SPLITT-OUT-X86-LSmitll_DFFT-IN X531-LSmitll_SPLITT-OUT-X86-LSmitll_DFFT-IN X86-LSmitll_DFFT-OUT-X114-LSmitll_SPLITT-INt LSmitll_DFFT

t902 X87-LSmitll_DFFT-OUT-X140-LSmitll_AND2T-INt 0 X87-LSmitll_DFFT-OUT-X140-LSmitll_AND2T-IN 0 z0=5 td=27.9ps
X87 X59-LSmitll_SPLITT-OUT-X87-LSmitll_DFFT-IN X459-LSmitll_SPLITT-OUT-X87-LSmitll_DFFT-IN X87-LSmitll_DFFT-OUT-X140-LSmitll_AND2T-INt LSmitll_DFFT

t903 X88-LSmitll_NOTT-OUT-X141-LSmitll_AND2T-INt 0 X88-LSmitll_NOTT-OUT-X141-LSmitll_AND2T-IN 0 z0=5 td=20.9ps
X88 X59-LSmitll_SPLITT-OUT-X88-LSmitll_NOTT-IN X460-LSmitll_SPLITT-OUT-X88-LSmitll_NOTT-IN X88-LSmitll_NOTT-OUT-X141-LSmitll_AND2T-INt LSmitll_NOTT

t904 X89-LSmitll_DFFT-OUT-X137-LSmitll_AND2T-INt 0 X89-LSmitll_DFFT-OUT-X137-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X89 X37-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-IN X313-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-IN X89-LSmitll_DFFT-OUT-X137-LSmitll_AND2T-INt LSmitll_DFFT

t905 X90-LSmitll_AND2T-OUT-X138-LSmitll_AND2T-INt 0 X90-LSmitll_AND2T-OUT-X138-LSmitll_AND2T-IN 0 z0=5 td=3.0ps
X90 X34-LSmitll_DFFT-OUT-X90-LSmitll_AND2T-IN X38-LSmitll_SPLITT-OUT-X90-LSmitll_AND2T-IN X350-LSmitll_SPLITT-OUT-X90-LSmitll_AND2T-IN X90-LSmitll_AND2T-OUT-X138-LSmitll_AND2T-INt LSmitll_AND2T

t906 X91-LSmitll_DFFT-OUT-X139-LSmitll_AND2T-INt 0 X91-LSmitll_DFFT-OUT-X139-LSmitll_AND2T-IN 0 z0=5 td=11.6ps
X91 X39-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-IN X314-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-IN X91-LSmitll_DFFT-OUT-X139-LSmitll_AND2T-INt LSmitll_DFFT

t907 X92-LSmitll_DFFT-OUT-X140-LSmitll_AND2T-INt 0 X92-LSmitll_DFFT-OUT-X140-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X92 X38-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-IN X343-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-IN X92-LSmitll_DFFT-OUT-X140-LSmitll_AND2T-INt LSmitll_DFFT

t908 X93-LSmitll_OR2T-OUT-X141-LSmitll_AND2T-INt 0 X93-LSmitll_OR2T-OUT-X141-LSmitll_AND2T-IN 0 z0=5 td=16.5ps
X93 X37-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-IN X39-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-IN X314-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-IN X93-LSmitll_OR2T-OUT-X141-LSmitll_AND2T-INt LSmitll_OR2T

t909 X94-LSmitll_SPLITT-OUT-X96-LSmitll_SPLITT-INt 0 X94-LSmitll_SPLITT-OUT-X96-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t910 X94-LSmitll_SPLITT-OUT-X95-LSmitll_SPLITT-INt 0 X94-LSmitll_SPLITT-OUT-X95-LSmitll_SPLITT-IN 0 z0=5 td=2.8ps
X94 X66-LSmitll_DFFT-OUT-X94-LSmitll_SPLITT-IN X94-LSmitll_SPLITT-OUT-X96-LSmitll_SPLITT-INt X94-LSmitll_SPLITT-OUT-X95-LSmitll_SPLITT-INt LSmitll_SPLITT

t911 X95-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-INt 0 X95-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-IN 0 z0=5 td=8.0ps
t912 X95-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-INt 0 X95-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-IN 0 z0=5 td=2.9ps
X95 X94-LSmitll_SPLITT-OUT-X95-LSmitll_SPLITT-IN X95-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-INt X95-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-INt LSmitll_SPLITT

t913 X96-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-INt 0 X96-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t914 X96-LSmitll_SPLITT-OUT-X125-LSmitll_AND2T-INt 0 X96-LSmitll_SPLITT-OUT-X125-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
X96 X94-LSmitll_SPLITT-OUT-X96-LSmitll_SPLITT-IN X96-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-INt X96-LSmitll_SPLITT-OUT-X125-LSmitll_AND2T-INt LSmitll_SPLITT

t915 X97-LSmitll_SPLITT-OUT-X238-LSmitll_OR2T-INt 0 X97-LSmitll_SPLITT-OUT-X238-LSmitll_OR2T-IN 0 z0=5 td=2.2ps
t916 X97-LSmitll_SPLITT-OUT-X98-LSmitll_SPLITT-INt 0 X97-LSmitll_SPLITT-OUT-X98-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X97 X67-LSmitll_DFFT-OUT-X97-LSmitll_SPLITT-IN X97-LSmitll_SPLITT-OUT-X238-LSmitll_OR2T-INt X97-LSmitll_SPLITT-OUT-X98-LSmitll_SPLITT-INt LSmitll_SPLITT

t917 X98-LSmitll_SPLITT-OUT-X134-LSmitll_AND2T-INt 0 X98-LSmitll_SPLITT-OUT-X134-LSmitll_AND2T-IN 0 z0=5 td=3.3ps
t918 X98-LSmitll_SPLITT-OUT-X131-LSmitll_AND2T-INt 0 X98-LSmitll_SPLITT-OUT-X131-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
X98 X97-LSmitll_SPLITT-OUT-X98-LSmitll_SPLITT-IN X98-LSmitll_SPLITT-OUT-X134-LSmitll_AND2T-INt X98-LSmitll_SPLITT-OUT-X131-LSmitll_AND2T-INt LSmitll_SPLITT

t919 X99-LSmitll_SPLITT-OUT-X101-LSmitll_SPLITT-INt 0 X99-LSmitll_SPLITT-OUT-X101-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t920 X99-LSmitll_SPLITT-OUT-X100-LSmitll_SPLITT-INt 0 X99-LSmitll_SPLITT-OUT-X100-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X99 X64-LSmitll_DFFT-OUT-X99-LSmitll_SPLITT-IN X99-LSmitll_SPLITT-OUT-X101-LSmitll_SPLITT-INt X99-LSmitll_SPLITT-OUT-X100-LSmitll_SPLITT-INt LSmitll_SPLITT

t921 X100-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-INt 0 X100-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-IN 0 z0=5 td=1.2ps
t922 X100-LSmitll_SPLITT-OUT-X116-LSmitll_DFFT-INt 0 X100-LSmitll_SPLITT-OUT-X116-LSmitll_DFFT-IN 0 z0=5 td=4.7ps
X100 X99-LSmitll_SPLITT-OUT-X100-LSmitll_SPLITT-IN X100-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-INt X100-LSmitll_SPLITT-OUT-X116-LSmitll_DFFT-INt LSmitll_SPLITT

t923 X101-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-INt 0 X101-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t924 X101-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt 0 X101-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN 0 z0=5 td=3.1ps
X101 X99-LSmitll_SPLITT-OUT-X101-LSmitll_SPLITT-IN X101-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-INt X101-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt LSmitll_SPLITT

t925 X102-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-INt 0 X102-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t926 X102-LSmitll_SPLITT-OUT-X103-LSmitll_SPLITT-INt 0 X102-LSmitll_SPLITT-OUT-X103-LSmitll_SPLITT-IN 0 z0=5 td=4.1ps
X102 X65-LSmitll_DFFT-OUT-X102-LSmitll_SPLITT-IN X102-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-INt X102-LSmitll_SPLITT-OUT-X103-LSmitll_SPLITT-INt LSmitll_SPLITT

t927 X103-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-INt 0 X103-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-IN 0 z0=5 td=3.3ps
t928 X103-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt 0 X103-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X103 X102-LSmitll_SPLITT-OUT-X103-LSmitll_SPLITT-IN X103-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-INt X103-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt LSmitll_SPLITT

t929 X104-LSmitll_SPLITT-OUT-X118-LSmitll_DFFT-INt 0 X104-LSmitll_SPLITT-OUT-X118-LSmitll_DFFT-IN 0 z0=5 td=2.5ps
t930 X104-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-INt 0 X104-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-IN 0 z0=5 td=4.8ps
X104 X60-LSmitll_DFFT-OUT-X104-LSmitll_SPLITT-IN X104-LSmitll_SPLITT-OUT-X118-LSmitll_DFFT-INt X104-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-INt LSmitll_SPLITT

t931 X105-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt 0 X105-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t932 X105-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt 0 X105-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
X105 X61-LSmitll_DFFT-OUT-X105-LSmitll_SPLITT-IN X105-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt X105-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt LSmitll_SPLITT

t933 X106-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt 0 X106-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN 0 z0=5 td=3.4ps
t934 X106-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-INt 0 X106-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-IN 0 z0=5 td=6.4ps
X106 X62-LSmitll_DFFT-OUT-X106-LSmitll_SPLITT-IN X106-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt X106-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-INt LSmitll_SPLITT

t935 X107-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-INt 0 X107-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
t936 X107-LSmitll_SPLITT-OUT-X108-LSmitll_SPLITT-INt 0 X107-LSmitll_SPLITT-OUT-X108-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X107 X63-LSmitll_DFFT-OUT-X107-LSmitll_SPLITT-IN X107-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-INt X107-LSmitll_SPLITT-OUT-X108-LSmitll_SPLITT-INt LSmitll_SPLITT

t937 X108-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt 0 X108-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN 0 z0=5 td=1.5ps
t938 X108-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-INt 0 X108-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
X108 X107-LSmitll_SPLITT-OUT-X108-LSmitll_SPLITT-IN X108-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt X108-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-INt LSmitll_SPLITT

t939 X109-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt 0 X109-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t940 X109-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-INt 0 X109-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-IN 0 z0=5 td=3.5ps
X109 X69-LSmitll_NOTT-OUT-X109-LSmitll_SPLITT-IN X109-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt X109-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-INt LSmitll_SPLITT

t941 X110-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt 0 X110-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
t942 X110-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-INt 0 X110-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
X110 X70-LSmitll_DFFT-OUT-X110-LSmitll_SPLITT-IN X110-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt X110-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-INt LSmitll_SPLITT

t943 X111-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt 0 X111-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN 0 z0=5 td=4.1ps
t944 X111-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-INt 0 X111-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X111 X74-LSmitll_DFFT-OUT-X111-LSmitll_SPLITT-IN X111-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt X111-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-INt LSmitll_SPLITT

t945 X112-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-INt 0 X112-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
t946 X112-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt 0 X112-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X112 X78-LSmitll_DFFT-OUT-X112-LSmitll_SPLITT-IN X112-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-INt X112-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt LSmitll_SPLITT

t947 X113-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt 0 X113-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN 0 z0=5 td=3.9ps
t948 X113-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-INt 0 X113-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-IN 0 z0=5 td=2.6ps
X113 X82-LSmitll_DFFT-OUT-X113-LSmitll_SPLITT-IN X113-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt X113-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-INt LSmitll_SPLITT

t949 X114-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-INt 0 X114-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-IN 0 z0=5 td=4.3ps
t950 X114-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt 0 X114-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN 0 z0=5 td=4.6ps
X114 X86-LSmitll_DFFT-OUT-X114-LSmitll_SPLITT-IN X114-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-INt X114-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt LSmitll_SPLITT

t951 X115-LSmitll_DFFT-OUT-X156-LSmitll_AND2T-INt 0 X115-LSmitll_DFFT-OUT-X156-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
X115 X68-LSmitll_DFFT-OUT-X115-LSmitll_DFFT-IN X400-LSmitll_SPLITT-OUT-X115-LSmitll_DFFT-IN X115-LSmitll_DFFT-OUT-X156-LSmitll_AND2T-INt LSmitll_DFFT

t952 X116-LSmitll_DFFT-OUT-X146-LSmitll_DFFT-INt 0 X116-LSmitll_DFFT-OUT-X146-LSmitll_DFFT-IN 0 z0=5 td=3.5ps
X116 X100-LSmitll_SPLITT-OUT-X116-LSmitll_DFFT-IN X551-LSmitll_SPLITT-OUT-X116-LSmitll_DFFT-IN X116-LSmitll_DFFT-OUT-X146-LSmitll_DFFT-INt LSmitll_DFFT


X117 X100-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-IN X104-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-IN X365-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-IN readt LSmitll_OR2T

t954 X118-LSmitll_DFFT-OUT-X147-LSmitll_DFFT-INt 0 X118-LSmitll_DFFT-OUT-X147-LSmitll_DFFT-IN 0 z0=5 td=3.3ps
X118 X104-LSmitll_SPLITT-OUT-X118-LSmitll_DFFT-IN X454-LSmitll_SPLITT-OUT-X118-LSmitll_DFFT-IN X118-LSmitll_DFFT-OUT-X147-LSmitll_DFFT-INt LSmitll_DFFT

t955 X119-LSmitll_AND2T-OUT-X149-LSmitll_DFFT-INt 0 X119-LSmitll_AND2T-OUT-X149-LSmitll_DFFT-IN 0 z0=5 td=4.6ps
X119 X95-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-IN X109-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-IN X363-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-IN X119-LSmitll_AND2T-OUT-X149-LSmitll_DFFT-INt LSmitll_AND2T

t956 X120-LSmitll_AND2T-OUT-X148-LSmitll_DFFT-INt 0 X120-LSmitll_AND2T-OUT-X148-LSmitll_DFFT-IN 0 z0=5 td=10.7ps
X120 X109-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN X105-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN X357-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN X120-LSmitll_AND2T-OUT-X148-LSmitll_DFFT-INt LSmitll_AND2T

t957 X121-LSmitll_AND2T-OUT-X151-LSmitll_DFFT-INt 0 X121-LSmitll_AND2T-OUT-X151-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X121 X95-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-IN X110-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-IN X473-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-IN X121-LSmitll_AND2T-OUT-X151-LSmitll_DFFT-INt LSmitll_AND2T

t958 X122-LSmitll_AND2T-OUT-X150-LSmitll_DFFT-INt 0 X122-LSmitll_AND2T-OUT-X150-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X122 X105-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN X110-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN X451-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN X122-LSmitll_AND2T-OUT-X150-LSmitll_DFFT-INt LSmitll_AND2T

t959 X123-LSmitll_AND2T-OUT-X152-LSmitll_OR2T-INt 0 X123-LSmitll_AND2T-OUT-X152-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X123 X106-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-IN X111-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-IN X334-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-IN X123-LSmitll_AND2T-OUT-X152-LSmitll_OR2T-INt LSmitll_AND2T

t960 X124-LSmitll_AND2T-OUT-X152-LSmitll_OR2T-INt 0 X124-LSmitll_AND2T-OUT-X152-LSmitll_OR2T-IN 0 z0=5 td=1.3ps
X124 X111-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN X101-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN X331-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN X124-LSmitll_AND2T-OUT-X152-LSmitll_OR2T-INt LSmitll_AND2T


X125 X73-LSmitll_DFFT-OUT-X125-LSmitll_AND2T-IN X96-LSmitll_SPLITT-OUT-X125-LSmitll_AND2T-IN X328-LSmitll_SPLITT-OUT-X125-LSmitll_AND2T-IN Imm0t LSmitll_AND2T

t962 X126-LSmitll_AND2T-OUT-X153-LSmitll_OR2T-INt 0 X126-LSmitll_AND2T-OUT-X153-LSmitll_OR2T-IN 0 z0=5 td=16.0ps
X126 X106-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN X112-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN X552-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN X126-LSmitll_AND2T-OUT-X153-LSmitll_OR2T-INt LSmitll_AND2T

t963 X127-LSmitll_AND2T-OUT-X153-LSmitll_OR2T-INt 0 X127-LSmitll_AND2T-OUT-X153-LSmitll_OR2T-IN 0 z0=5 td=1.3ps
X127 X101-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-IN X112-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-IN X337-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-IN X127-LSmitll_AND2T-OUT-X153-LSmitll_OR2T-INt LSmitll_AND2T


X128 X77-LSmitll_DFFT-OUT-X128-LSmitll_AND2T-IN X96-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-IN X365-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-IN Imm1t LSmitll_AND2T

t965 X129-LSmitll_AND2T-OUT-X154-LSmitll_OR2T-INt 0 X129-LSmitll_AND2T-OUT-X154-LSmitll_OR2T-IN 0 z0=5 td=13.9ps
X129 X108-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-IN X113-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-IN X404-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-IN X129-LSmitll_AND2T-OUT-X154-LSmitll_OR2T-INt LSmitll_AND2T

t966 X130-LSmitll_AND2T-OUT-X154-LSmitll_OR2T-INt 0 X130-LSmitll_AND2T-OUT-X154-LSmitll_OR2T-IN 0 z0=5 td=16.5ps
X130 X113-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN X103-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN X502-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN X130-LSmitll_AND2T-OUT-X154-LSmitll_OR2T-INt LSmitll_AND2T


X131 X81-LSmitll_DFFT-OUT-X131-LSmitll_AND2T-IN X98-LSmitll_SPLITT-OUT-X131-LSmitll_AND2T-IN X508-LSmitll_SPLITT-OUT-X131-LSmitll_AND2T-IN Imm2t LSmitll_AND2T

t968 X132-LSmitll_AND2T-OUT-X155-LSmitll_OR2T-INt 0 X132-LSmitll_AND2T-OUT-X155-LSmitll_OR2T-IN 0 z0=5 td=7.5ps
X132 X108-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN X114-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN X508-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN X132-LSmitll_AND2T-OUT-X155-LSmitll_OR2T-INt LSmitll_AND2T

t969 X133-LSmitll_AND2T-OUT-X155-LSmitll_OR2T-INt 0 X133-LSmitll_AND2T-OUT-X155-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X133 X103-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-IN X114-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-IN X509-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-IN X133-LSmitll_AND2T-OUT-X155-LSmitll_OR2T-INt LSmitll_AND2T


X134 X85-LSmitll_DFFT-OUT-X134-LSmitll_AND2T-IN X98-LSmitll_SPLITT-OUT-X134-LSmitll_AND2T-IN X531-LSmitll_SPLITT-OUT-X134-LSmitll_AND2T-IN Imm3t LSmitll_AND2T

t971 X135-LSmitll_OR2T-OUT-X156-LSmitll_AND2T-INt 0 X135-LSmitll_OR2T-OUT-X156-LSmitll_AND2T-IN 0 z0=5 td=3.9ps
X135 X71-LSmitll_DFFT-OUT-X135-LSmitll_OR2T-IN X75-LSmitll_DFFT-OUT-X135-LSmitll_OR2T-IN X378-LSmitll_SPLITT-OUT-X135-LSmitll_OR2T-IN X135-LSmitll_OR2T-OUT-X156-LSmitll_AND2T-INt LSmitll_OR2T

t972 X136-LSmitll_DFFT-OUT-X157-LSmitll_OR2T-INt 0 X136-LSmitll_DFFT-OUT-X157-LSmitll_OR2T-IN 0 z0=5 td=5.0ps
X136 X79-LSmitll_DFFT-OUT-X136-LSmitll_DFFT-IN X317-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-IN X136-LSmitll_DFFT-OUT-X157-LSmitll_OR2T-INt LSmitll_DFFT

t973 X137-LSmitll_AND2T-OUT-X157-LSmitll_OR2T-INt 0 X137-LSmitll_AND2T-OUT-X157-LSmitll_OR2T-IN 0 z0=5 td=8.6ps
X137 X80-LSmitll_NOTT-OUT-X137-LSmitll_AND2T-IN X89-LSmitll_DFFT-OUT-X137-LSmitll_AND2T-IN X313-LSmitll_SPLITT-OUT-X137-LSmitll_AND2T-IN X137-LSmitll_AND2T-OUT-X157-LSmitll_OR2T-INt LSmitll_AND2T

t974 X138-LSmitll_AND2T-OUT-X158-LSmitll_OR2T-INt 0 X138-LSmitll_AND2T-OUT-X158-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X138 X83-LSmitll_DFFT-OUT-X138-LSmitll_AND2T-IN X90-LSmitll_AND2T-OUT-X138-LSmitll_AND2T-IN X430-LSmitll_SPLITT-OUT-X138-LSmitll_AND2T-IN X138-LSmitll_AND2T-OUT-X158-LSmitll_OR2T-INt LSmitll_AND2T

t975 X139-LSmitll_AND2T-OUT-X158-LSmitll_OR2T-INt 0 X139-LSmitll_AND2T-OUT-X158-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X139 X84-LSmitll_NOTT-OUT-X139-LSmitll_AND2T-IN X91-LSmitll_DFFT-OUT-X139-LSmitll_AND2T-IN X343-LSmitll_SPLITT-OUT-X139-LSmitll_AND2T-IN X139-LSmitll_AND2T-OUT-X158-LSmitll_OR2T-INt LSmitll_AND2T

t976 X140-LSmitll_AND2T-OUT-X159-LSmitll_OR2T-INt 0 X140-LSmitll_AND2T-OUT-X159-LSmitll_OR2T-IN 0 z0=5 td=0.9ps
X140 X87-LSmitll_DFFT-OUT-X140-LSmitll_AND2T-IN X92-LSmitll_DFFT-OUT-X140-LSmitll_AND2T-IN X342-LSmitll_SPLITT-OUT-X140-LSmitll_AND2T-IN X140-LSmitll_AND2T-OUT-X159-LSmitll_OR2T-INt LSmitll_AND2T

t977 X141-LSmitll_AND2T-OUT-X159-LSmitll_OR2T-INt 0 X141-LSmitll_AND2T-OUT-X159-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X141 X88-LSmitll_NOTT-OUT-X141-LSmitll_AND2T-IN X93-LSmitll_OR2T-OUT-X141-LSmitll_AND2T-IN X321-LSmitll_SPLITT-OUT-X141-LSmitll_AND2T-IN X141-LSmitll_AND2T-OUT-X159-LSmitll_OR2T-INt LSmitll_AND2T

t978 X142-LSmitll_DFFT-OUT-X160-LSmitll_DFFT-INt 0 X142-LSmitll_DFFT-OUT-X160-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X142 X72-LSmitll_DFFT-OUT-X142-LSmitll_DFFT-IN X401-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-IN X142-LSmitll_DFFT-OUT-X160-LSmitll_DFFT-INt LSmitll_DFFT

t979 X143-LSmitll_DFFT-OUT-X161-LSmitll_DFFT-INt 0 X143-LSmitll_DFFT-OUT-X161-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X143 X76-LSmitll_DFFT-OUT-X143-LSmitll_DFFT-IN X378-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-IN X143-LSmitll_DFFT-OUT-X161-LSmitll_DFFT-INt LSmitll_DFFT

t980 X144-LSmitll_DFFT-OUT-X220-LSmitll_DFFT-INt 0 X144-LSmitll_DFFT-OUT-X220-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X144 X107-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-IN X393-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-IN X144-LSmitll_DFFT-OUT-X220-LSmitll_DFFT-INt LSmitll_DFFT

t981 X145-LSmitll_DFFT-OUT-X162-LSmitll_DFFT-INt 0 X145-LSmitll_DFFT-OUT-X162-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X145 X102-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-IN X553-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-IN X145-LSmitll_DFFT-OUT-X162-LSmitll_DFFT-INt LSmitll_DFFT

t982 X146-LSmitll_DFFT-OUT-X164-LSmitll_DFFT-INt 0 X146-LSmitll_DFFT-OUT-X164-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X146 X116-LSmitll_DFFT-OUT-X146-LSmitll_DFFT-IN X489-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-IN X146-LSmitll_DFFT-OUT-X164-LSmitll_DFFT-INt LSmitll_DFFT

t983 X147-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-INt 0 X147-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-IN 0 z0=5 td=3.4ps
X147 X118-LSmitll_DFFT-OUT-X147-LSmitll_DFFT-IN X489-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-IN X147-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-INt LSmitll_DFFT

t984 X148-LSmitll_DFFT-OUT-X166-LSmitll_DFFT-INt 0 X148-LSmitll_DFFT-OUT-X166-LSmitll_DFFT-IN 0 z0=5 td=4.7ps
X148 X120-LSmitll_AND2T-OUT-X148-LSmitll_DFFT-IN X335-LSmitll_SPLITT-OUT-X148-LSmitll_DFFT-IN X148-LSmitll_DFFT-OUT-X166-LSmitll_DFFT-INt LSmitll_DFFT

t985 X149-LSmitll_DFFT-OUT-X167-LSmitll_DFFT-INt 0 X149-LSmitll_DFFT-OUT-X167-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X149 X119-LSmitll_AND2T-OUT-X149-LSmitll_DFFT-IN X352-LSmitll_SPLITT-OUT-X149-LSmitll_DFFT-IN X149-LSmitll_DFFT-OUT-X167-LSmitll_DFFT-INt LSmitll_DFFT

t986 X150-LSmitll_DFFT-OUT-X168-LSmitll_DFFT-INt 0 X150-LSmitll_DFFT-OUT-X168-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X150 X122-LSmitll_AND2T-OUT-X150-LSmitll_DFFT-IN X448-LSmitll_SPLITT-OUT-X150-LSmitll_DFFT-IN X150-LSmitll_DFFT-OUT-X168-LSmitll_DFFT-INt LSmitll_DFFT

t987 X151-LSmitll_DFFT-OUT-X169-LSmitll_DFFT-INt 0 X151-LSmitll_DFFT-OUT-X169-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X151 X121-LSmitll_AND2T-OUT-X151-LSmitll_DFFT-IN X474-LSmitll_SPLITT-OUT-X151-LSmitll_DFFT-IN X151-LSmitll_DFFT-OUT-X169-LSmitll_DFFT-INt LSmitll_DFFT

t988 X152-LSmitll_OR2T-OUT-X170-LSmitll_DFFT-INt 0 X152-LSmitll_OR2T-OUT-X170-LSmitll_DFFT-IN 0 z0=5 td=2.4ps
X152 X123-LSmitll_AND2T-OUT-X152-LSmitll_OR2T-IN X124-LSmitll_AND2T-OUT-X152-LSmitll_OR2T-IN X330-LSmitll_SPLITT-OUT-X152-LSmitll_OR2T-IN X152-LSmitll_OR2T-OUT-X170-LSmitll_DFFT-INt LSmitll_OR2T

t989 X153-LSmitll_OR2T-OUT-X171-LSmitll_DFFT-INt 0 X153-LSmitll_OR2T-OUT-X171-LSmitll_DFFT-IN 0 z0=5 td=4.6ps
X153 X126-LSmitll_AND2T-OUT-X153-LSmitll_OR2T-IN X127-LSmitll_AND2T-OUT-X153-LSmitll_OR2T-IN X331-LSmitll_SPLITT-OUT-X153-LSmitll_OR2T-IN X153-LSmitll_OR2T-OUT-X171-LSmitll_DFFT-INt LSmitll_OR2T

t990 X154-LSmitll_OR2T-OUT-X172-LSmitll_DFFT-INt 0 X154-LSmitll_OR2T-OUT-X172-LSmitll_DFFT-IN 0 z0=5 td=10.5ps
X154 X129-LSmitll_AND2T-OUT-X154-LSmitll_OR2T-IN X130-LSmitll_AND2T-OUT-X154-LSmitll_OR2T-IN X509-LSmitll_SPLITT-OUT-X154-LSmitll_OR2T-IN X154-LSmitll_OR2T-OUT-X172-LSmitll_DFFT-INt LSmitll_OR2T

t991 X155-LSmitll_OR2T-OUT-X163-LSmitll_SPLITT-INt 0 X155-LSmitll_OR2T-OUT-X163-LSmitll_SPLITT-IN 0 z0=5 td=7.0ps
X155 X132-LSmitll_AND2T-OUT-X155-LSmitll_OR2T-IN X133-LSmitll_AND2T-OUT-X155-LSmitll_OR2T-IN X519-LSmitll_SPLITT-OUT-X155-LSmitll_OR2T-IN X155-LSmitll_OR2T-OUT-X163-LSmitll_SPLITT-INt LSmitll_OR2T

t992 X156-LSmitll_AND2T-OUT-X175-LSmitll_DFFT-INt 0 X156-LSmitll_AND2T-OUT-X175-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
X156 X115-LSmitll_DFFT-OUT-X156-LSmitll_AND2T-IN X135-LSmitll_OR2T-OUT-X156-LSmitll_AND2T-IN X379-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-IN X156-LSmitll_AND2T-OUT-X175-LSmitll_DFFT-INt LSmitll_AND2T

t993 X157-LSmitll_OR2T-OUT-X177-LSmitll_DFFT-INt 0 X157-LSmitll_OR2T-OUT-X177-LSmitll_DFFT-IN 0 z0=5 td=3.4ps
X157 X136-LSmitll_DFFT-OUT-X157-LSmitll_OR2T-IN X137-LSmitll_AND2T-OUT-X157-LSmitll_OR2T-IN X321-LSmitll_SPLITT-OUT-X157-LSmitll_OR2T-IN X157-LSmitll_OR2T-OUT-X177-LSmitll_DFFT-INt LSmitll_OR2T

t994 X158-LSmitll_OR2T-OUT-X176-LSmitll_OR2T-INt 0 X158-LSmitll_OR2T-OUT-X176-LSmitll_OR2T-IN 0 z0=5 td=3.5ps
X158 X138-LSmitll_AND2T-OUT-X158-LSmitll_OR2T-IN X139-LSmitll_AND2T-OUT-X158-LSmitll_OR2T-IN X349-LSmitll_SPLITT-OUT-X158-LSmitll_OR2T-IN X158-LSmitll_OR2T-OUT-X176-LSmitll_OR2T-INt LSmitll_OR2T

t995 X159-LSmitll_OR2T-OUT-X176-LSmitll_OR2T-INt 0 X159-LSmitll_OR2T-OUT-X176-LSmitll_OR2T-IN 0 z0=5 td=7.9ps
X159 X140-LSmitll_AND2T-OUT-X159-LSmitll_OR2T-IN X141-LSmitll_AND2T-OUT-X159-LSmitll_OR2T-IN X342-LSmitll_SPLITT-OUT-X159-LSmitll_OR2T-IN X159-LSmitll_OR2T-OUT-X176-LSmitll_OR2T-INt LSmitll_OR2T

t996 X160-LSmitll_DFFT-OUT-X178-LSmitll_DFFT-INt 0 X160-LSmitll_DFFT-OUT-X178-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X160 X142-LSmitll_DFFT-OUT-X160-LSmitll_DFFT-IN X404-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-IN X160-LSmitll_DFFT-OUT-X178-LSmitll_DFFT-INt LSmitll_DFFT

t997 X161-LSmitll_DFFT-OUT-X179-LSmitll_DFFT-INt 0 X161-LSmitll_DFFT-OUT-X179-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X161 X143-LSmitll_DFFT-OUT-X161-LSmitll_DFFT-IN X372-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-IN X161-LSmitll_DFFT-OUT-X179-LSmitll_DFFT-INt LSmitll_DFFT

t998 X162-LSmitll_DFFT-OUT-X206-LSmitll_DFFT-INt 0 X162-LSmitll_DFFT-OUT-X206-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X162 X145-LSmitll_DFFT-OUT-X162-LSmitll_DFFT-IN X519-LSmitll_SPLITT-OUT-X162-LSmitll_DFFT-IN X162-LSmitll_DFFT-OUT-X206-LSmitll_DFFT-INt LSmitll_DFFT

t999 X163-LSmitll_SPLITT-OUT-X174-LSmitll_DFFT-INt 0 X163-LSmitll_SPLITT-OUT-X174-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
t1000 X163-LSmitll_SPLITT-OUT-X173-LSmitll_DFFT-INt 0 X163-LSmitll_SPLITT-OUT-X173-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X163 X155-LSmitll_OR2T-OUT-X163-LSmitll_SPLITT-IN X163-LSmitll_SPLITT-OUT-X174-LSmitll_DFFT-INt X163-LSmitll_SPLITT-OUT-X173-LSmitll_DFFT-INt LSmitll_SPLITT

t1001 X164-LSmitll_DFFT-OUT-X181-LSmitll_DFFT-INt 0 X164-LSmitll_DFFT-OUT-X181-LSmitll_DFFT-IN 0 z0=5 td=5.3ps
X164 X146-LSmitll_DFFT-OUT-X164-LSmitll_DFFT-IN X488-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-IN X164-LSmitll_DFFT-OUT-X181-LSmitll_DFFT-INt LSmitll_DFFT

t1002 X165-LSmitll_DFFT-OUT-X182-LSmitll_DFFT-INt 0 X165-LSmitll_DFFT-OUT-X182-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X165 X147-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-IN X495-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-IN X165-LSmitll_DFFT-OUT-X182-LSmitll_DFFT-INt LSmitll_DFFT

t1003 X166-LSmitll_DFFT-OUT-X183-LSmitll_DFFT-INt 0 X166-LSmitll_DFFT-OUT-X183-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X166 X148-LSmitll_DFFT-OUT-X166-LSmitll_DFFT-IN X323-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-IN X166-LSmitll_DFFT-OUT-X183-LSmitll_DFFT-INt LSmitll_DFFT

t1004 X167-LSmitll_DFFT-OUT-X311-LSmitll_OR2T-INt 0 X167-LSmitll_DFFT-OUT-X311-LSmitll_OR2T-IN 0 z0=5 td=25.3ps
X167 X149-LSmitll_DFFT-OUT-X167-LSmitll_DFFT-IN X346-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-IN X167-LSmitll_DFFT-OUT-X311-LSmitll_OR2T-INt LSmitll_DFFT

t1005 X168-LSmitll_DFFT-OUT-X184-LSmitll_DFFT-INt 0 X168-LSmitll_DFFT-OUT-X184-LSmitll_DFFT-IN 0 z0=5 td=3.8ps
X168 X150-LSmitll_DFFT-OUT-X168-LSmitll_DFFT-IN X447-LSmitll_SPLITT-OUT-X168-LSmitll_DFFT-IN X168-LSmitll_DFFT-OUT-X184-LSmitll_DFFT-INt LSmitll_DFFT

t1006 X169-LSmitll_DFFT-OUT-X312-LSmitll_OR2T-INt 0 X169-LSmitll_DFFT-OUT-X312-LSmitll_OR2T-IN 0 z0=5 td=3.7ps
X169 X151-LSmitll_DFFT-OUT-X169-LSmitll_DFFT-IN X479-LSmitll_SPLITT-OUT-X169-LSmitll_DFFT-IN X169-LSmitll_DFFT-OUT-X312-LSmitll_OR2T-INt LSmitll_DFFT

t1007 X170-LSmitll_DFFT-OUT-X185-LSmitll_DFFT-INt 0 X170-LSmitll_DFFT-OUT-X185-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X170 X152-LSmitll_OR2T-OUT-X170-LSmitll_DFFT-IN X328-LSmitll_SPLITT-OUT-X170-LSmitll_DFFT-IN X170-LSmitll_DFFT-OUT-X185-LSmitll_DFFT-INt LSmitll_DFFT

t1008 X171-LSmitll_DFFT-OUT-X186-LSmitll_DFFT-INt 0 X171-LSmitll_DFFT-OUT-X186-LSmitll_DFFT-IN 0 z0=5 td=2.7ps
X171 X153-LSmitll_OR2T-OUT-X171-LSmitll_DFFT-IN X371-LSmitll_SPLITT-OUT-X171-LSmitll_DFFT-IN X171-LSmitll_DFFT-OUT-X186-LSmitll_DFFT-INt LSmitll_DFFT

t1009 X172-LSmitll_DFFT-OUT-X187-LSmitll_DFFT-INt 0 X172-LSmitll_DFFT-OUT-X187-LSmitll_DFFT-IN 0 z0=5 td=2.4ps
X172 X154-LSmitll_OR2T-OUT-X172-LSmitll_DFFT-IN X539-LSmitll_SPLITT-OUT-X172-LSmitll_DFFT-IN X172-LSmitll_DFFT-OUT-X187-LSmitll_DFFT-INt LSmitll_DFFT

t1010 X173-LSmitll_DFFT-OUT-X180-LSmitll_SPLITT-INt 0 X173-LSmitll_DFFT-OUT-X180-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X173 X163-LSmitll_SPLITT-OUT-X173-LSmitll_DFFT-IN X533-LSmitll_SPLITT-OUT-X173-LSmitll_DFFT-IN X173-LSmitll_DFFT-OUT-X180-LSmitll_SPLITT-INt LSmitll_DFFT

t1011 X174-LSmitll_DFFT-OUT-X190-LSmitll_DFFT-INt 0 X174-LSmitll_DFFT-OUT-X190-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X174 X163-LSmitll_SPLITT-OUT-X174-LSmitll_DFFT-IN X533-LSmitll_SPLITT-OUT-X174-LSmitll_DFFT-IN X174-LSmitll_DFFT-OUT-X190-LSmitll_DFFT-INt LSmitll_DFFT

t1012 X175-LSmitll_DFFT-OUT-X191-LSmitll_DFFT-INt 0 X175-LSmitll_DFFT-OUT-X191-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X175 X156-LSmitll_AND2T-OUT-X175-LSmitll_DFFT-IN X554-LSmitll_SPLITT-OUT-X175-LSmitll_DFFT-IN X175-LSmitll_DFFT-OUT-X191-LSmitll_DFFT-INt LSmitll_DFFT

t1013 X176-LSmitll_OR2T-OUT-X192-LSmitll_OR2T-INt 0 X176-LSmitll_OR2T-OUT-X192-LSmitll_OR2T-IN 0 z0=5 td=3.9ps
X176 X158-LSmitll_OR2T-OUT-X176-LSmitll_OR2T-IN X159-LSmitll_OR2T-OUT-X176-LSmitll_OR2T-IN X352-LSmitll_SPLITT-OUT-X176-LSmitll_OR2T-IN X176-LSmitll_OR2T-OUT-X192-LSmitll_OR2T-INt LSmitll_OR2T

t1014 X177-LSmitll_DFFT-OUT-X192-LSmitll_OR2T-INt 0 X177-LSmitll_DFFT-OUT-X192-LSmitll_OR2T-IN 0 z0=5 td=2.3ps
X177 X157-LSmitll_OR2T-OUT-X177-LSmitll_DFFT-IN X345-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-IN X177-LSmitll_DFFT-OUT-X192-LSmitll_OR2T-INt LSmitll_DFFT

t1015 X178-LSmitll_DFFT-OUT-X193-LSmitll_DFFT-INt 0 X178-LSmitll_DFFT-OUT-X193-LSmitll_DFFT-IN 0 z0=5 td=15.0ps
X178 X160-LSmitll_DFFT-OUT-X178-LSmitll_DFFT-IN X407-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-IN X178-LSmitll_DFFT-OUT-X193-LSmitll_DFFT-INt LSmitll_DFFT

t1016 X179-LSmitll_DFFT-OUT-X194-LSmitll_DFFT-INt 0 X179-LSmitll_DFFT-OUT-X194-LSmitll_DFFT-IN 0 z0=5 td=14.8ps
X179 X161-LSmitll_DFFT-OUT-X179-LSmitll_DFFT-IN X372-LSmitll_SPLITT-OUT-X179-LSmitll_DFFT-IN X179-LSmitll_DFFT-OUT-X194-LSmitll_DFFT-INt LSmitll_DFFT

t1017 X180-LSmitll_SPLITT-OUT-X189-LSmitll_DFFT-INt 0 X180-LSmitll_SPLITT-OUT-X189-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
t1018 X180-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-INt 0 X180-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X180 X173-LSmitll_DFFT-OUT-X180-LSmitll_SPLITT-IN X180-LSmitll_SPLITT-OUT-X189-LSmitll_DFFT-INt X180-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-INt LSmitll_SPLITT

t1019 X181-LSmitll_DFFT-OUT-X197-LSmitll_DFFT-INt 0 X181-LSmitll_DFFT-OUT-X197-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X181 X164-LSmitll_DFFT-OUT-X181-LSmitll_DFFT-IN X408-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-IN X181-LSmitll_DFFT-OUT-X197-LSmitll_DFFT-INt LSmitll_DFFT

t1020 X182-LSmitll_DFFT-OUT-X198-LSmitll_DFFT-INt 0 X182-LSmitll_DFFT-OUT-X198-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X182 X165-LSmitll_DFFT-OUT-X182-LSmitll_DFFT-IN X555-LSmitll_SPLITT-OUT-X182-LSmitll_DFFT-IN X182-LSmitll_DFFT-OUT-X198-LSmitll_DFFT-INt LSmitll_DFFT

t1021 X183-LSmitll_DFFT-OUT-X199-LSmitll_DFFT-INt 0 X183-LSmitll_DFFT-OUT-X199-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X183 X166-LSmitll_DFFT-OUT-X183-LSmitll_DFFT-IN X317-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-IN X183-LSmitll_DFFT-OUT-X199-LSmitll_DFFT-INt LSmitll_DFFT

t1022 X184-LSmitll_DFFT-OUT-X200-LSmitll_DFFT-INt 0 X184-LSmitll_DFFT-OUT-X200-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X184 X168-LSmitll_DFFT-OUT-X184-LSmitll_DFFT-IN X444-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-IN X184-LSmitll_DFFT-OUT-X200-LSmitll_DFFT-INt LSmitll_DFFT


X185 X170-LSmitll_DFFT-OUT-X185-LSmitll_DFFT-IN X327-LSmitll_SPLITT-OUT-X185-LSmitll_DFFT-IN Op_Aritht LSmitll_DFFT


X186 X171-LSmitll_DFFT-OUT-X186-LSmitll_DFFT-IN X371-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-IN Op_Andt LSmitll_DFFT


X187 X172-LSmitll_DFFT-OUT-X187-LSmitll_DFFT-IN X556-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-IN Op_Xort LSmitll_DFFT


X188 X180-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-IN X539-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-IN Cmpl_b0t LSmitll_DFFT


X189 X180-LSmitll_SPLITT-OUT-X189-LSmitll_DFFT-IN X511-LSmitll_SPLITT-OUT-X189-LSmitll_DFFT-IN Cmpl_b1t LSmitll_DFFT


X190 X174-LSmitll_DFFT-OUT-X190-LSmitll_DFFT-IN X557-LSmitll_SPLITT-OUT-X190-LSmitll_DFFT-IN Cint LSmitll_DFFT

t1029 X191-LSmitll_DFFT-OUT-X196-LSmitll_SPLITT-INt 0 X191-LSmitll_DFFT-OUT-X196-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X191 X175-LSmitll_DFFT-OUT-X191-LSmitll_DFFT-IN X381-LSmitll_SPLITT-OUT-X191-LSmitll_DFFT-IN X191-LSmitll_DFFT-OUT-X196-LSmitll_SPLITT-INt LSmitll_DFFT

t1030 X192-LSmitll_OR2T-OUT-X195-LSmitll_SPLITT-INt 0 X192-LSmitll_OR2T-OUT-X195-LSmitll_SPLITT-IN 0 z0=5 td=12.7ps
X192 X176-LSmitll_OR2T-OUT-X192-LSmitll_OR2T-IN X177-LSmitll_DFFT-OUT-X192-LSmitll_OR2T-IN X346-LSmitll_SPLITT-OUT-X192-LSmitll_OR2T-IN X192-LSmitll_OR2T-OUT-X195-LSmitll_SPLITT-INt LSmitll_OR2T

t1031 X193-LSmitll_DFFT-OUT-X204-LSmitll_DFFT-INt 0 X193-LSmitll_DFFT-OUT-X204-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X193 X178-LSmitll_DFFT-OUT-X193-LSmitll_DFFT-IN X498-LSmitll_SPLITT-OUT-X193-LSmitll_DFFT-IN X193-LSmitll_DFFT-OUT-X204-LSmitll_DFFT-INt LSmitll_DFFT

t1032 X194-LSmitll_DFFT-OUT-X205-LSmitll_DFFT-INt 0 X194-LSmitll_DFFT-OUT-X205-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X194 X179-LSmitll_DFFT-OUT-X194-LSmitll_DFFT-IN X374-LSmitll_SPLITT-OUT-X194-LSmitll_DFFT-IN X194-LSmitll_DFFT-OUT-X205-LSmitll_DFFT-INt LSmitll_DFFT

t1033 X195-LSmitll_SPLITT-OUT-X203-LSmitll_NOTT-INt 0 X195-LSmitll_SPLITT-OUT-X203-LSmitll_NOTT-IN 0 z0=5 td=1.7ps
t1034 X195-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-INt 0 X195-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-IN 0 z0=5 td=2.9ps
X195 X192-LSmitll_OR2T-OUT-X195-LSmitll_SPLITT-IN X195-LSmitll_SPLITT-OUT-X203-LSmitll_NOTT-INt X195-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-INt LSmitll_SPLITT

t1035 X196-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-INt 0 X196-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-IN 0 z0=5 td=3.3ps
t1036 X196-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-INt 0 X196-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X196 X191-LSmitll_DFFT-OUT-X196-LSmitll_SPLITT-IN X196-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-INt X196-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-INt LSmitll_SPLITT

t1037 X197-LSmitll_DFFT-OUT-X210-LSmitll_DFFT-INt 0 X197-LSmitll_DFFT-OUT-X210-LSmitll_DFFT-IN 0 z0=5 td=3.5ps
X197 X181-LSmitll_DFFT-OUT-X197-LSmitll_DFFT-IN X408-LSmitll_SPLITT-OUT-X197-LSmitll_DFFT-IN X197-LSmitll_DFFT-OUT-X210-LSmitll_DFFT-INt LSmitll_DFFT

t1038 X198-LSmitll_DFFT-OUT-X211-LSmitll_DFFT-INt 0 X198-LSmitll_DFFT-OUT-X211-LSmitll_DFFT-IN 0 z0=5 td=4.9ps
X198 X182-LSmitll_DFFT-OUT-X198-LSmitll_DFFT-IN X516-LSmitll_SPLITT-OUT-X198-LSmitll_DFFT-IN X198-LSmitll_DFFT-OUT-X211-LSmitll_DFFT-INt LSmitll_DFFT

t1039 X199-LSmitll_DFFT-OUT-X212-LSmitll_DFFT-INt 0 X199-LSmitll_DFFT-OUT-X212-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X199 X183-LSmitll_DFFT-OUT-X199-LSmitll_DFFT-IN X316-LSmitll_SPLITT-OUT-X199-LSmitll_DFFT-IN X199-LSmitll_DFFT-OUT-X212-LSmitll_DFFT-INt LSmitll_DFFT

t1040 X200-LSmitll_DFFT-OUT-X213-LSmitll_DFFT-INt 0 X200-LSmitll_DFFT-OUT-X213-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
X200 X184-LSmitll_DFFT-OUT-X200-LSmitll_DFFT-IN X444-LSmitll_SPLITT-OUT-X200-LSmitll_DFFT-IN X200-LSmitll_DFFT-OUT-X213-LSmitll_DFFT-INt LSmitll_DFFT

t1041 X201-LSmitll_DFFT-OUT-X208-LSmitll_SPLITT-INt 0 X201-LSmitll_DFFT-OUT-X208-LSmitll_SPLITT-IN 0 z0=5 td=4.4ps
X201 X196-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-IN X403-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-IN X201-LSmitll_DFFT-OUT-X208-LSmitll_SPLITT-INt LSmitll_DFFT

t1042 X202-LSmitll_AND2T-OUT-X207-LSmitll_SPLITT-INt 0 X202-LSmitll_AND2T-OUT-X207-LSmitll_SPLITT-IN 0 z0=5 td=5.6ps
X202 X196-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-IN X195-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-IN X403-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-IN X202-LSmitll_AND2T-OUT-X207-LSmitll_SPLITT-INt LSmitll_AND2T

t1043 X203-LSmitll_NOTT-OUT-X214-LSmitll_AND2T-INt 0 X203-LSmitll_NOTT-OUT-X214-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
X203 X195-LSmitll_SPLITT-OUT-X203-LSmitll_NOTT-IN X410-LSmitll_SPLITT-OUT-X203-LSmitll_NOTT-IN X203-LSmitll_NOTT-OUT-X214-LSmitll_AND2T-INt LSmitll_NOTT

t1044 X204-LSmitll_DFFT-OUT-X218-LSmitll_AND2T-INt 0 X204-LSmitll_DFFT-OUT-X218-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X204 X193-LSmitll_DFFT-OUT-X204-LSmitll_DFFT-IN X492-LSmitll_SPLITT-OUT-X204-LSmitll_DFFT-IN X204-LSmitll_DFFT-OUT-X218-LSmitll_AND2T-INt LSmitll_DFFT

t1045 X205-LSmitll_DFFT-OUT-X219-LSmitll_AND2T-INt 0 X205-LSmitll_DFFT-OUT-X219-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
X205 X194-LSmitll_DFFT-OUT-X205-LSmitll_DFFT-IN X374-LSmitll_SPLITT-OUT-X205-LSmitll_DFFT-IN X205-LSmitll_DFFT-OUT-X219-LSmitll_AND2T-INt LSmitll_DFFT

t1046 X206-LSmitll_DFFT-OUT-X221-LSmitll_DFFT-INt 0 X206-LSmitll_DFFT-OUT-X221-LSmitll_DFFT-IN 0 z0=5 td=5.2ps
X206 X162-LSmitll_DFFT-OUT-X206-LSmitll_DFFT-IN X520-LSmitll_SPLITT-OUT-X206-LSmitll_DFFT-IN X206-LSmitll_DFFT-OUT-X221-LSmitll_DFFT-INt LSmitll_DFFT

t1047 X207-LSmitll_SPLITT-OUT-X215-LSmitll_DFFT-INt 0 X207-LSmitll_SPLITT-OUT-X215-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
t1048 X207-LSmitll_SPLITT-OUT-X209-LSmitll_SPLITT-INt 0 X207-LSmitll_SPLITT-OUT-X209-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X207 X202-LSmitll_AND2T-OUT-X207-LSmitll_SPLITT-IN X207-LSmitll_SPLITT-OUT-X215-LSmitll_DFFT-INt X207-LSmitll_SPLITT-OUT-X209-LSmitll_SPLITT-INt LSmitll_SPLITT

t1049 X208-LSmitll_SPLITT-OUT-X217-LSmitll_DFFT-INt 0 X208-LSmitll_SPLITT-OUT-X217-LSmitll_DFFT-IN 0 z0=5 td=3.2ps
t1050 X208-LSmitll_SPLITT-OUT-X214-LSmitll_AND2T-INt 0 X208-LSmitll_SPLITT-OUT-X214-LSmitll_AND2T-IN 0 z0=5 td=1.1ps
X208 X201-LSmitll_DFFT-OUT-X208-LSmitll_SPLITT-IN X208-LSmitll_SPLITT-OUT-X217-LSmitll_DFFT-INt X208-LSmitll_SPLITT-OUT-X214-LSmitll_AND2T-INt LSmitll_SPLITT

t1051 X209-LSmitll_SPLITT-OUT-X219-LSmitll_AND2T-INt 0 X209-LSmitll_SPLITT-OUT-X219-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1052 X209-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-INt 0 X209-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
X209 X207-LSmitll_SPLITT-OUT-X209-LSmitll_SPLITT-IN X209-LSmitll_SPLITT-OUT-X219-LSmitll_AND2T-INt X209-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-INt LSmitll_SPLITT

t1053 X210-LSmitll_DFFT-OUT-X222-LSmitll_DFFT-INt 0 X210-LSmitll_DFFT-OUT-X222-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X210 X197-LSmitll_DFFT-OUT-X210-LSmitll_DFFT-IN X488-LSmitll_SPLITT-OUT-X210-LSmitll_DFFT-IN X210-LSmitll_DFFT-OUT-X222-LSmitll_DFFT-INt LSmitll_DFFT

t1054 X211-LSmitll_DFFT-OUT-X223-LSmitll_DFFT-INt 0 X211-LSmitll_DFFT-OUT-X223-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X211 X198-LSmitll_DFFT-OUT-X211-LSmitll_DFFT-IN X523-LSmitll_SPLITT-OUT-X211-LSmitll_DFFT-IN X211-LSmitll_DFFT-OUT-X223-LSmitll_DFFT-INt LSmitll_DFFT

t1055 X212-LSmitll_DFFT-OUT-X224-LSmitll_DFFT-INt 0 X212-LSmitll_DFFT-OUT-X224-LSmitll_DFFT-IN 0 z0=5 td=6.5ps
X212 X199-LSmitll_DFFT-OUT-X212-LSmitll_DFFT-IN X327-LSmitll_SPLITT-OUT-X212-LSmitll_DFFT-IN X212-LSmitll_DFFT-OUT-X224-LSmitll_DFFT-INt LSmitll_DFFT

t1056 X213-LSmitll_DFFT-OUT-X225-LSmitll_DFFT-INt 0 X213-LSmitll_DFFT-OUT-X225-LSmitll_DFFT-IN 0 z0=5 td=5.5ps
X213 X200-LSmitll_DFFT-OUT-X213-LSmitll_DFFT-IN X363-LSmitll_SPLITT-OUT-X213-LSmitll_DFFT-IN X213-LSmitll_DFFT-OUT-X225-LSmitll_DFFT-INt LSmitll_DFFT

t1057 X214-LSmitll_AND2T-OUT-X230-LSmitll_OR2T-INt 0 X214-LSmitll_AND2T-OUT-X230-LSmitll_OR2T-IN 0 z0=5 td=5.1ps
X214 X203-LSmitll_NOTT-OUT-X214-LSmitll_AND2T-IN X208-LSmitll_SPLITT-OUT-X214-LSmitll_AND2T-IN X410-LSmitll_SPLITT-OUT-X214-LSmitll_AND2T-IN X214-LSmitll_AND2T-OUT-X230-LSmitll_OR2T-INt LSmitll_AND2T

t1058 X215-LSmitll_DFFT-OUT-X228-LSmitll_DFFT-INt 0 X215-LSmitll_DFFT-OUT-X228-LSmitll_DFFT-IN 0 z0=5 td=3.1ps
X215 X207-LSmitll_SPLITT-OUT-X215-LSmitll_DFFT-IN X386-LSmitll_SPLITT-OUT-X215-LSmitll_DFFT-IN X215-LSmitll_DFFT-OUT-X228-LSmitll_DFFT-INt LSmitll_DFFT

t1059 X216-LSmitll_OR2T-OUT-X229-LSmitll_AND2T-INt 0 X216-LSmitll_OR2T-OUT-X229-LSmitll_AND2T-IN 0 z0=5 td=5.6ps
X216 X295-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-IN X296-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-IN X420-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-IN X216-LSmitll_OR2T-OUT-X229-LSmitll_AND2T-INt LSmitll_OR2T

t1060 X217-LSmitll_DFFT-OUT-X229-LSmitll_AND2T-INt 0 X217-LSmitll_DFFT-OUT-X229-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X217 X208-LSmitll_SPLITT-OUT-X217-LSmitll_DFFT-IN X415-LSmitll_SPLITT-OUT-X217-LSmitll_DFFT-IN X217-LSmitll_DFFT-OUT-X229-LSmitll_AND2T-INt LSmitll_DFFT

t1061 X218-LSmitll_AND2T-OUT-X230-LSmitll_OR2T-INt 0 X218-LSmitll_AND2T-OUT-X230-LSmitll_OR2T-IN 0 z0=5 td=21.5ps
X218 X204-LSmitll_DFFT-OUT-X218-LSmitll_AND2T-IN X209-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-IN X491-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-IN X218-LSmitll_AND2T-OUT-X230-LSmitll_OR2T-INt LSmitll_AND2T

t1062 X219-LSmitll_AND2T-OUT-X231-LSmitll_DFFT-INt 0 X219-LSmitll_AND2T-OUT-X231-LSmitll_DFFT-IN 0 z0=5 td=5.2ps
X219 X205-LSmitll_DFFT-OUT-X219-LSmitll_AND2T-IN X209-LSmitll_SPLITT-OUT-X219-LSmitll_AND2T-IN X375-LSmitll_SPLITT-OUT-X219-LSmitll_AND2T-IN X219-LSmitll_AND2T-OUT-X231-LSmitll_DFFT-INt LSmitll_AND2T

t1063 X220-LSmitll_DFFT-OUT-X233-LSmitll_OR2T-INt 0 X220-LSmitll_DFFT-OUT-X233-LSmitll_OR2T-IN 0 z0=5 td=0.9ps
X220 X144-LSmitll_DFFT-OUT-X220-LSmitll_DFFT-IN X381-LSmitll_SPLITT-OUT-X220-LSmitll_DFFT-IN X220-LSmitll_DFFT-OUT-X233-LSmitll_OR2T-INt LSmitll_DFFT

t1064 X221-LSmitll_DFFT-OUT-X226-LSmitll_DFFT-INt 0 X221-LSmitll_DFFT-OUT-X226-LSmitll_DFFT-IN 0 z0=5 td=33.4ps
X221 X206-LSmitll_DFFT-OUT-X221-LSmitll_DFFT-IN X498-LSmitll_SPLITT-OUT-X221-LSmitll_DFFT-IN X221-LSmitll_DFFT-OUT-X226-LSmitll_DFFT-INt LSmitll_DFFT

t1065 X222-LSmitll_DFFT-OUT-X234-LSmitll_DFFT-INt 0 X222-LSmitll_DFFT-OUT-X234-LSmitll_DFFT-IN 0 z0=5 td=13.9ps
X222 X210-LSmitll_DFFT-OUT-X222-LSmitll_DFFT-IN X491-LSmitll_SPLITT-OUT-X222-LSmitll_DFFT-IN X222-LSmitll_DFFT-OUT-X234-LSmitll_DFFT-INt LSmitll_DFFT

t1066 X223-LSmitll_DFFT-OUT-X235-LSmitll_DFFT-INt 0 X223-LSmitll_DFFT-OUT-X235-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X223 X211-LSmitll_DFFT-OUT-X223-LSmitll_DFFT-IN X517-LSmitll_SPLITT-OUT-X223-LSmitll_DFFT-IN X223-LSmitll_DFFT-OUT-X235-LSmitll_DFFT-INt LSmitll_DFFT

t1067 X224-LSmitll_DFFT-OUT-X236-LSmitll_DFFT-INt 0 X224-LSmitll_DFFT-OUT-X236-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X224 X212-LSmitll_DFFT-OUT-X224-LSmitll_DFFT-IN X323-LSmitll_SPLITT-OUT-X224-LSmitll_DFFT-IN X224-LSmitll_DFFT-OUT-X236-LSmitll_DFFT-INt LSmitll_DFFT

t1068 X225-LSmitll_DFFT-OUT-X237-LSmitll_DFFT-INt 0 X225-LSmitll_DFFT-OUT-X237-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X225 X213-LSmitll_DFFT-OUT-X225-LSmitll_DFFT-IN X445-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-IN X225-LSmitll_DFFT-OUT-X237-LSmitll_DFFT-INt LSmitll_DFFT

t1069 X226-LSmitll_DFFT-OUT-X227-LSmitll_DFFT-INt 0 X226-LSmitll_DFFT-OUT-X227-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X226 X221-LSmitll_DFFT-OUT-X226-LSmitll_DFFT-IN X385-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-IN X226-LSmitll_DFFT-OUT-X227-LSmitll_DFFT-INt LSmitll_DFFT

t1070 X227-LSmitll_DFFT-OUT-X233-LSmitll_OR2T-INt 0 X227-LSmitll_DFFT-OUT-X233-LSmitll_OR2T-IN 0 z0=5 td=3.9ps
X227 X226-LSmitll_DFFT-OUT-X227-LSmitll_DFFT-IN X386-LSmitll_SPLITT-OUT-X227-LSmitll_DFFT-IN X227-LSmitll_DFFT-OUT-X233-LSmitll_OR2T-INt LSmitll_DFFT

t1071 X228-LSmitll_DFFT-OUT-X240-LSmitll_OR2T-INt 0 X228-LSmitll_DFFT-OUT-X240-LSmitll_OR2T-IN 0 z0=5 td=5.1ps
X228 X215-LSmitll_DFFT-OUT-X228-LSmitll_DFFT-IN X389-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-IN X228-LSmitll_DFFT-OUT-X240-LSmitll_OR2T-INt LSmitll_DFFT

t1072 X229-LSmitll_AND2T-OUT-X240-LSmitll_OR2T-INt 0 X229-LSmitll_AND2T-OUT-X240-LSmitll_OR2T-IN 0 z0=5 td=1.3ps
X229 X216-LSmitll_OR2T-OUT-X229-LSmitll_AND2T-IN X217-LSmitll_DFFT-OUT-X229-LSmitll_AND2T-IN X414-LSmitll_SPLITT-OUT-X229-LSmitll_AND2T-IN X229-LSmitll_AND2T-OUT-X240-LSmitll_OR2T-INt LSmitll_AND2T

t1073 X230-LSmitll_OR2T-OUT-X241-LSmitll_OR2T-INt 0 X230-LSmitll_OR2T-OUT-X241-LSmitll_OR2T-IN 0 z0=5 td=15.0ps
X230 X214-LSmitll_AND2T-OUT-X230-LSmitll_OR2T-IN X218-LSmitll_AND2T-OUT-X230-LSmitll_OR2T-IN X420-LSmitll_SPLITT-OUT-X230-LSmitll_OR2T-IN X230-LSmitll_OR2T-OUT-X241-LSmitll_OR2T-INt LSmitll_OR2T

t1074 X231-LSmitll_DFFT-OUT-X242-LSmitll_DFFT-INt 0 X231-LSmitll_DFFT-OUT-X242-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X231 X219-LSmitll_AND2T-OUT-X231-LSmitll_DFFT-IN X388-LSmitll_SPLITT-OUT-X231-LSmitll_DFFT-IN X231-LSmitll_DFFT-OUT-X242-LSmitll_DFFT-INt LSmitll_DFFT

t1075 X232-LSmitll_OR2T-OUT-X243-LSmitll_AND2T-INt 0 X232-LSmitll_OR2T-OUT-X243-LSmitll_AND2T-IN 0 z0=5 td=2.7ps
X232 X295-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-IN X296-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-IN X421-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-IN X232-LSmitll_OR2T-OUT-X243-LSmitll_AND2T-INt LSmitll_OR2T

t1076 X233-LSmitll_OR2T-OUT-X238-LSmitll_OR2T-INt 0 X233-LSmitll_OR2T-OUT-X238-LSmitll_OR2T-IN 0 z0=5 td=17.0ps
X233 X220-LSmitll_DFFT-OUT-X233-LSmitll_OR2T-IN X227-LSmitll_DFFT-OUT-X233-LSmitll_OR2T-IN X375-LSmitll_SPLITT-OUT-X233-LSmitll_OR2T-IN X233-LSmitll_OR2T-OUT-X238-LSmitll_OR2T-INt LSmitll_OR2T

t1077 X234-LSmitll_DFFT-OUT-X246-LSmitll_DFFT-INt 0 X234-LSmitll_DFFT-OUT-X246-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X234 X222-LSmitll_DFFT-OUT-X234-LSmitll_DFFT-IN X520-LSmitll_SPLITT-OUT-X234-LSmitll_DFFT-IN X234-LSmitll_DFFT-OUT-X246-LSmitll_DFFT-INt LSmitll_DFFT

t1078 X235-LSmitll_DFFT-OUT-X247-LSmitll_DFFT-INt 0 X235-LSmitll_DFFT-OUT-X247-LSmitll_DFFT-IN 0 z0=5 td=6.8ps
X235 X223-LSmitll_DFFT-OUT-X235-LSmitll_DFFT-IN X476-LSmitll_SPLITT-OUT-X235-LSmitll_DFFT-IN X235-LSmitll_DFFT-OUT-X247-LSmitll_DFFT-INt LSmitll_DFFT

t1079 X236-LSmitll_DFFT-OUT-X248-LSmitll_DFFT-INt 0 X236-LSmitll_DFFT-OUT-X248-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X236 X224-LSmitll_DFFT-OUT-X236-LSmitll_DFFT-IN X558-LSmitll_SPLITT-OUT-X236-LSmitll_DFFT-IN X236-LSmitll_DFFT-OUT-X248-LSmitll_DFFT-INt LSmitll_DFFT

t1080 X237-LSmitll_DFFT-OUT-X249-LSmitll_DFFT-INt 0 X237-LSmitll_DFFT-OUT-X249-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X237 X225-LSmitll_DFFT-OUT-X237-LSmitll_DFFT-IN X445-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-IN X237-LSmitll_DFFT-OUT-X249-LSmitll_DFFT-INt LSmitll_DFFT

t1081 X238-LSmitll_OR2T-OUT-X239-LSmitll_SPLITT-INt 0 X238-LSmitll_OR2T-OUT-X239-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X238 X97-LSmitll_SPLITT-OUT-X238-LSmitll_OR2T-IN X233-LSmitll_OR2T-OUT-X238-LSmitll_OR2T-IN X502-LSmitll_SPLITT-OUT-X238-LSmitll_OR2T-IN X238-LSmitll_OR2T-OUT-X239-LSmitll_SPLITT-INt LSmitll_OR2T

t1082 X239-LSmitll_SPLITT-OUT-X243-LSmitll_AND2T-INt 0 X239-LSmitll_SPLITT-OUT-X243-LSmitll_AND2T-IN 0 z0=5 td=2.9ps
t1083 X239-LSmitll_SPLITT-OUT-X241-LSmitll_OR2T-INt 0 X239-LSmitll_SPLITT-OUT-X241-LSmitll_OR2T-IN 0 z0=5 td=1.4ps
X239 X238-LSmitll_OR2T-OUT-X239-LSmitll_SPLITT-IN X239-LSmitll_SPLITT-OUT-X243-LSmitll_AND2T-INt X239-LSmitll_SPLITT-OUT-X241-LSmitll_OR2T-INt LSmitll_SPLITT

t1084 X240-LSmitll_OR2T-OUT-X253-LSmitll_OR2T-INt 0 X240-LSmitll_OR2T-OUT-X253-LSmitll_OR2T-IN 0 z0=5 td=1.3ps
X240 X228-LSmitll_DFFT-OUT-X240-LSmitll_OR2T-IN X229-LSmitll_AND2T-OUT-X240-LSmitll_OR2T-IN X393-LSmitll_SPLITT-OUT-X240-LSmitll_OR2T-IN X240-LSmitll_OR2T-OUT-X253-LSmitll_OR2T-INt LSmitll_OR2T

t1085 X241-LSmitll_OR2T-OUT-X245-LSmitll_SPLITT-INt 0 X241-LSmitll_OR2T-OUT-X245-LSmitll_SPLITT-IN 0 z0=5 td=13.4ps
X241 X230-LSmitll_OR2T-OUT-X241-LSmitll_OR2T-IN X239-LSmitll_SPLITT-OUT-X241-LSmitll_OR2T-IN X421-LSmitll_SPLITT-OUT-X241-LSmitll_OR2T-IN X241-LSmitll_OR2T-OUT-X245-LSmitll_SPLITT-INt LSmitll_OR2T

t1086 X242-LSmitll_DFFT-OUT-X252-LSmitll_XORT-INt 0 X242-LSmitll_DFFT-OUT-X252-LSmitll_XORT-IN 0 z0=5 td=17.0ps
X242 X231-LSmitll_DFFT-OUT-X242-LSmitll_DFFT-IN X385-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-IN X242-LSmitll_DFFT-OUT-X252-LSmitll_XORT-INt LSmitll_DFFT

t1087 X243-LSmitll_AND2T-OUT-X253-LSmitll_OR2T-INt 0 X243-LSmitll_AND2T-OUT-X253-LSmitll_OR2T-IN 0 z0=5 td=15.1ps
X243 X232-LSmitll_OR2T-OUT-X243-LSmitll_AND2T-IN X239-LSmitll_SPLITT-OUT-X243-LSmitll_AND2T-IN X415-LSmitll_SPLITT-OUT-X243-LSmitll_AND2T-IN X243-LSmitll_AND2T-OUT-X253-LSmitll_OR2T-INt LSmitll_AND2T

t1088 X244-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-INt 0 X244-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1089 X244-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-INt 0 X244-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-IN 0 z0=5 td=3.6ps
X244 X291-LSmitll_DFFT-OUT-X244-LSmitll_SPLITT-IN X244-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-INt X244-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-INt LSmitll_SPLITT

t1090 X245-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-INt 0 X245-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-IN 0 z0=5 td=3.6ps
t1091 X245-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-INt 0 X245-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-IN 0 z0=5 td=2.1ps
X245 X241-LSmitll_OR2T-OUT-X245-LSmitll_SPLITT-IN X245-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-INt X245-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-INt LSmitll_SPLITT

t1092 X246-LSmitll_DFFT-OUT-X254-LSmitll_DFFT-INt 0 X246-LSmitll_DFFT-OUT-X254-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X246 X234-LSmitll_DFFT-OUT-X246-LSmitll_DFFT-IN X526-LSmitll_SPLITT-OUT-X246-LSmitll_DFFT-IN X246-LSmitll_DFFT-OUT-X254-LSmitll_DFFT-INt LSmitll_DFFT

t1093 X247-LSmitll_DFFT-OUT-X255-LSmitll_DFFT-INt 0 X247-LSmitll_DFFT-OUT-X255-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X247 X235-LSmitll_DFFT-OUT-X247-LSmitll_DFFT-IN X516-LSmitll_SPLITT-OUT-X247-LSmitll_DFFT-IN X247-LSmitll_DFFT-OUT-X255-LSmitll_DFFT-INt LSmitll_DFFT

t1094 X248-LSmitll_DFFT-OUT-X256-LSmitll_DFFT-INt 0 X248-LSmitll_DFFT-OUT-X256-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X248 X236-LSmitll_DFFT-OUT-X248-LSmitll_DFFT-IN X356-LSmitll_SPLITT-OUT-X248-LSmitll_DFFT-IN X248-LSmitll_DFFT-OUT-X256-LSmitll_DFFT-INt LSmitll_DFFT

t1095 X249-LSmitll_DFFT-OUT-X257-LSmitll_DFFT-INt 0 X249-LSmitll_DFFT-OUT-X257-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X249 X237-LSmitll_DFFT-OUT-X249-LSmitll_DFFT-IN X440-LSmitll_SPLITT-OUT-X249-LSmitll_DFFT-IN X249-LSmitll_DFFT-OUT-X257-LSmitll_DFFT-INt LSmitll_DFFT

t1096 X250-LSmitll_XORT-OUT-X260-LSmitll_DFFT-INt 0 X250-LSmitll_XORT-OUT-X260-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X250 X244-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-IN X245-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-IN X559-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-IN X250-LSmitll_XORT-OUT-X260-LSmitll_DFFT-INt LSmitll_XORT

t1097 X251-LSmitll_AND2T-OUT-X259-LSmitll_XORT-INt 0 X251-LSmitll_AND2T-OUT-X259-LSmitll_XORT-IN 0 z0=5 td=17.7ps
X251 X244-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-IN X245-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-IN X530-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-IN X251-LSmitll_AND2T-OUT-X259-LSmitll_XORT-INt LSmitll_AND2T

t1098 X252-LSmitll_XORT-OUT-X259-LSmitll_XORT-INt 0 X252-LSmitll_XORT-OUT-X259-LSmitll_XORT-IN 0 z0=5 td=2.5ps
X252 X242-LSmitll_DFFT-OUT-X252-LSmitll_XORT-IN X292-LSmitll_DFFT-OUT-X252-LSmitll_XORT-IN X414-LSmitll_SPLITT-OUT-X252-LSmitll_XORT-IN X252-LSmitll_XORT-OUT-X259-LSmitll_XORT-INt LSmitll_XORT

t1099 X253-LSmitll_OR2T-OUT-X258-LSmitll_SPLITT-INt 0 X253-LSmitll_OR2T-OUT-X258-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X253 X240-LSmitll_OR2T-OUT-X253-LSmitll_OR2T-IN X243-LSmitll_AND2T-OUT-X253-LSmitll_OR2T-IN X392-LSmitll_SPLITT-OUT-X253-LSmitll_OR2T-IN X253-LSmitll_OR2T-OUT-X258-LSmitll_SPLITT-INt LSmitll_OR2T

t1100 X254-LSmitll_DFFT-OUT-X269-LSmitll_DFFT-INt 0 X254-LSmitll_DFFT-OUT-X269-LSmitll_DFFT-IN 0 z0=5 td=14.9ps
X254 X246-LSmitll_DFFT-OUT-X254-LSmitll_DFFT-IN X526-LSmitll_SPLITT-OUT-X254-LSmitll_DFFT-IN X254-LSmitll_DFFT-OUT-X269-LSmitll_DFFT-INt LSmitll_DFFT

t1101 X255-LSmitll_DFFT-OUT-X270-LSmitll_DFFT-INt 0 X255-LSmitll_DFFT-OUT-X270-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X255 X247-LSmitll_DFFT-OUT-X255-LSmitll_DFFT-IN X496-LSmitll_SPLITT-OUT-X255-LSmitll_DFFT-IN X255-LSmitll_DFFT-OUT-X270-LSmitll_DFFT-INt LSmitll_DFFT

t1102 X256-LSmitll_DFFT-OUT-X271-LSmitll_DFFT-INt 0 X256-LSmitll_DFFT-OUT-X271-LSmitll_DFFT-IN 0 z0=5 td=14.5ps
X256 X248-LSmitll_DFFT-OUT-X256-LSmitll_DFFT-IN X356-LSmitll_SPLITT-OUT-X256-LSmitll_DFFT-IN X256-LSmitll_DFFT-OUT-X271-LSmitll_DFFT-INt LSmitll_DFFT

t1103 X257-LSmitll_DFFT-OUT-X272-LSmitll_DFFT-INt 0 X257-LSmitll_DFFT-OUT-X272-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X257 X249-LSmitll_DFFT-OUT-X257-LSmitll_DFFT-IN X452-LSmitll_SPLITT-OUT-X257-LSmitll_DFFT-IN X257-LSmitll_DFFT-OUT-X272-LSmitll_DFFT-INt LSmitll_DFFT

t1104 X258-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-INt 0 X258-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
t1105 X258-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-INt 0 X258-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
X258 X253-LSmitll_OR2T-OUT-X258-LSmitll_SPLITT-IN X258-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-INt X258-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-INt LSmitll_SPLITT

t1106 X259-LSmitll_XORT-OUT-X266-LSmitll_SPLITT-INt 0 X259-LSmitll_XORT-OUT-X266-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X259 X251-LSmitll_AND2T-OUT-X259-LSmitll_XORT-IN X252-LSmitll_XORT-OUT-X259-LSmitll_XORT-IN X417-LSmitll_SPLITT-OUT-X259-LSmitll_XORT-IN X259-LSmitll_XORT-OUT-X266-LSmitll_SPLITT-INt LSmitll_XORT

t1107 X260-LSmitll_DFFT-OUT-X265-LSmitll_SPLITT-INt 0 X260-LSmitll_DFFT-OUT-X265-LSmitll_SPLITT-IN 0 z0=5 td=10.0ps
X260 X250-LSmitll_XORT-OUT-X260-LSmitll_DFFT-IN X537-LSmitll_SPLITT-OUT-X260-LSmitll_DFFT-IN X260-LSmitll_DFFT-OUT-X265-LSmitll_SPLITT-INt LSmitll_DFFT

t1108 X261-LSmitll_DFFT-OUT-X263-LSmitll_SPLITT-INt 0 X261-LSmitll_DFFT-OUT-X263-LSmitll_SPLITT-IN 0 z0=5 td=3.4ps
X261 X258-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-IN X560-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-IN X261-LSmitll_DFFT-OUT-X263-LSmitll_SPLITT-INt LSmitll_DFFT

t1109 X262-LSmitll_DFFT-OUT-X264-LSmitll_SPLITT-INt 0 X262-LSmitll_DFFT-OUT-X264-LSmitll_SPLITT-IN 0 z0=5 td=6.2ps
X262 X258-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-IN X388-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-IN X262-LSmitll_DFFT-OUT-X264-LSmitll_SPLITT-INt LSmitll_DFFT

t1110 X263-LSmitll_SPLITT-OUT-X279-LSmitll_SPLITT-INt 0 X263-LSmitll_SPLITT-OUT-X279-LSmitll_SPLITT-IN 0 z0=5 td=3.6ps
t1111 X263-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-INt 0 X263-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X263 X261-LSmitll_DFFT-OUT-X263-LSmitll_SPLITT-IN X263-LSmitll_SPLITT-OUT-X279-LSmitll_SPLITT-INt X263-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-INt LSmitll_SPLITT

t1112 X264-LSmitll_SPLITT-OUT-X282-LSmitll_SPLITT-INt 0 X264-LSmitll_SPLITT-OUT-X282-LSmitll_SPLITT-IN 0 z0=5 td=6.3ps
t1113 X264-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-INt 0 X264-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X264 X262-LSmitll_DFFT-OUT-X264-LSmitll_SPLITT-IN X264-LSmitll_SPLITT-OUT-X282-LSmitll_SPLITT-INt X264-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-INt LSmitll_SPLITT

t1114 X265-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-INt 0 X265-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1115 X265-LSmitll_SPLITT-OUT-X267-LSmitll_SPLITT-INt 0 X265-LSmitll_SPLITT-OUT-X267-LSmitll_SPLITT-IN 0 z0=5 td=5.5ps
X265 X260-LSmitll_DFFT-OUT-X265-LSmitll_SPLITT-IN X265-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-INt X265-LSmitll_SPLITT-OUT-X267-LSmitll_SPLITT-INt LSmitll_SPLITT

t1116 X266-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-INt 0 X266-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1117 X266-LSmitll_SPLITT-OUT-X268-LSmitll_SPLITT-INt 0 X266-LSmitll_SPLITT-OUT-X268-LSmitll_SPLITT-IN 0 z0=5 td=5.3ps
X266 X259-LSmitll_XORT-OUT-X266-LSmitll_SPLITT-IN X266-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-INt X266-LSmitll_SPLITT-OUT-X268-LSmitll_SPLITT-INt LSmitll_SPLITT

t1118 X267-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-INt 0 X267-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t1119 X267-LSmitll_SPLITT-OUT-X273-LSmitll_DFFT-INt 0 X267-LSmitll_SPLITT-OUT-X273-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X267 X265-LSmitll_SPLITT-OUT-X267-LSmitll_SPLITT-IN X267-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-INt X267-LSmitll_SPLITT-OUT-X273-LSmitll_DFFT-INt LSmitll_SPLITT

t1120 X268-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-INt 0 X268-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
t1121 X268-LSmitll_SPLITT-OUT-X275-LSmitll_DFFT-INt 0 X268-LSmitll_SPLITT-OUT-X275-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X268 X266-LSmitll_SPLITT-OUT-X268-LSmitll_SPLITT-IN X268-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-INt X268-LSmitll_SPLITT-OUT-X275-LSmitll_DFFT-INt LSmitll_SPLITT

t1122 X269-LSmitll_DFFT-OUT-X285-LSmitll_DFFT-INt 0 X269-LSmitll_DFFT-OUT-X285-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X269 X254-LSmitll_DFFT-OUT-X269-LSmitll_DFFT-IN X536-LSmitll_SPLITT-OUT-X269-LSmitll_DFFT-IN X269-LSmitll_DFFT-OUT-X285-LSmitll_DFFT-INt LSmitll_DFFT

t1123 X270-LSmitll_DFFT-OUT-X286-LSmitll_DFFT-INt 0 X270-LSmitll_DFFT-OUT-X286-LSmitll_DFFT-IN 0 z0=5 td=4.9ps
X270 X255-LSmitll_DFFT-OUT-X270-LSmitll_DFFT-IN X496-LSmitll_SPLITT-OUT-X270-LSmitll_DFFT-IN X270-LSmitll_DFFT-OUT-X286-LSmitll_DFFT-INt LSmitll_DFFT

t1124 X271-LSmitll_DFFT-OUT-X287-LSmitll_DFFT-INt 0 X271-LSmitll_DFFT-OUT-X287-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X271 X256-LSmitll_DFFT-OUT-X271-LSmitll_DFFT-IN X440-LSmitll_SPLITT-OUT-X271-LSmitll_DFFT-IN X271-LSmitll_DFFT-OUT-X287-LSmitll_DFFT-INt LSmitll_DFFT

t1125 X272-LSmitll_DFFT-OUT-X288-LSmitll_DFFT-INt 0 X272-LSmitll_DFFT-OUT-X288-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X272 X257-LSmitll_DFFT-OUT-X272-LSmitll_DFFT-IN X473-LSmitll_SPLITT-OUT-X272-LSmitll_DFFT-IN X272-LSmitll_DFFT-OUT-X288-LSmitll_DFFT-INt LSmitll_DFFT


X273 X267-LSmitll_SPLITT-OUT-X273-LSmitll_DFFT-IN X423-LSmitll_SPLITT-OUT-X273-LSmitll_DFFT-IN nextInstrAddr0_0t LSmitll_DFFT


X274 X267-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-IN X505-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-IN nextInstrAddr0_1t LSmitll_DFFT


X275 X268-LSmitll_SPLITT-OUT-X275-LSmitll_DFFT-IN X423-LSmitll_SPLITT-OUT-X275-LSmitll_DFFT-IN nextInstrAddr1_0t LSmitll_DFFT


X276 X268-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-IN X395-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-IN nextInstrAddr1_1t LSmitll_DFFT


X277 X263-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-IN X417-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-IN readNextInstr0t LSmitll_DFFT


X278 X264-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-IN X389-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-IN readNextInstr1t LSmitll_DFFT

t1132 X279-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-INt 0 X279-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1133 X279-LSmitll_SPLITT-OUT-X280-LSmitll_NDROT-INt 0 X279-LSmitll_SPLITT-OUT-X280-LSmitll_NDROT-IN 0 z0=5 td=5.4ps
X279 X263-LSmitll_SPLITT-OUT-X279-LSmitll_SPLITT-IN X279-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-INt X279-LSmitll_SPLITT-OUT-X280-LSmitll_NDROT-INt LSmitll_SPLITT

t1134 X280-LSmitll_NDROT-OUT-X289-LSmitll_SPLITT-INt 0 X280-LSmitll_NDROT-OUT-X289-LSmitll_SPLITT-IN 0 z0=5 td=4.0ps
X280 X281-LSmitll_AND2T-OUT-X280-LSmitll_NDROT-IN X279-LSmitll_SPLITT-OUT-X280-LSmitll_NDROT-IN X503-LSmitll_SPLITT-OUT-X280-LSmitll_NDROT-IN X280-LSmitll_NDROT-OUT-X289-LSmitll_SPLITT-INt LSmitll_NDROT

t1135 X281-LSmitll_AND2T-OUT-X280-LSmitll_NDROT-INt 0 X281-LSmitll_AND2T-OUT-X280-LSmitll_NDROT-IN 0 z0=5 td=3.6ps
X281 X265-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-IN X279-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-IN X505-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-IN X281-LSmitll_AND2T-OUT-X280-LSmitll_NDROT-INt LSmitll_AND2T

t1136 X282-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-INt 0 X282-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-IN 0 z0=5 td=4.9ps
t1137 X282-LSmitll_SPLITT-OUT-X283-LSmitll_NDROT-INt 0 X282-LSmitll_SPLITT-OUT-X283-LSmitll_NDROT-IN 0 z0=5 td=3.6ps
X282 X264-LSmitll_SPLITT-OUT-X282-LSmitll_SPLITT-IN X282-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-INt X282-LSmitll_SPLITT-OUT-X283-LSmitll_NDROT-INt LSmitll_SPLITT

t1138 X283-LSmitll_NDROT-OUT-X290-LSmitll_SPLITT-INt 0 X283-LSmitll_NDROT-OUT-X290-LSmitll_SPLITT-IN 0 z0=5 td=10.3ps
X283 X284-LSmitll_AND2T-OUT-X283-LSmitll_NDROT-IN X282-LSmitll_SPLITT-OUT-X283-LSmitll_NDROT-IN X392-LSmitll_SPLITT-OUT-X283-LSmitll_NDROT-IN X283-LSmitll_NDROT-OUT-X290-LSmitll_SPLITT-INt LSmitll_NDROT

t1139 X284-LSmitll_AND2T-OUT-X283-LSmitll_NDROT-INt 0 X284-LSmitll_AND2T-OUT-X283-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
X284 X266-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-IN X282-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-IN X395-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-IN X284-LSmitll_AND2T-OUT-X283-LSmitll_NDROT-INt LSmitll_AND2T

t1140 X285-LSmitll_DFFT-OUT-X297-LSmitll_DFFT-INt 0 X285-LSmitll_DFFT-OUT-X297-LSmitll_DFFT-IN 0 z0=5 td=4.2ps
X285 X269-LSmitll_DFFT-OUT-X285-LSmitll_DFFT-IN X561-LSmitll_SPLITT-OUT-X285-LSmitll_DFFT-IN X285-LSmitll_DFFT-OUT-X297-LSmitll_DFFT-INt LSmitll_DFFT

t1141 X286-LSmitll_DFFT-OUT-X298-LSmitll_DFFT-INt 0 X286-LSmitll_DFFT-OUT-X298-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X286 X270-LSmitll_DFFT-OUT-X286-LSmitll_DFFT-IN X517-LSmitll_SPLITT-OUT-X286-LSmitll_DFFT-IN X286-LSmitll_DFFT-OUT-X298-LSmitll_DFFT-INt LSmitll_DFFT

t1142 X287-LSmitll_DFFT-OUT-X299-LSmitll_DFFT-INt 0 X287-LSmitll_DFFT-OUT-X299-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X287 X271-LSmitll_DFFT-OUT-X287-LSmitll_DFFT-IN X562-LSmitll_SPLITT-OUT-X287-LSmitll_DFFT-IN X287-LSmitll_DFFT-OUT-X299-LSmitll_DFFT-INt LSmitll_DFFT

t1143 X288-LSmitll_DFFT-OUT-X300-LSmitll_DFFT-INt 0 X288-LSmitll_DFFT-OUT-X300-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X288 X272-LSmitll_DFFT-OUT-X288-LSmitll_DFFT-IN X463-LSmitll_SPLITT-OUT-X288-LSmitll_DFFT-IN X288-LSmitll_DFFT-OUT-X300-LSmitll_DFFT-INt LSmitll_DFFT

t1144 X289-LSmitll_SPLITT-OUT-X293-LSmitll_NOTT-INt 0 X289-LSmitll_SPLITT-OUT-X293-LSmitll_NOTT-IN 0 z0=5 td=1.2ps
t1145 X289-LSmitll_SPLITT-OUT-X291-LSmitll_DFFT-INt 0 X289-LSmitll_SPLITT-OUT-X291-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X289 X280-LSmitll_NDROT-OUT-X289-LSmitll_SPLITT-IN X289-LSmitll_SPLITT-OUT-X293-LSmitll_NOTT-INt X289-LSmitll_SPLITT-OUT-X291-LSmitll_DFFT-INt LSmitll_SPLITT

t1146 X290-LSmitll_SPLITT-OUT-X294-LSmitll_NOTT-INt 0 X290-LSmitll_SPLITT-OUT-X294-LSmitll_NOTT-IN 0 z0=5 td=5.2ps
t1147 X290-LSmitll_SPLITT-OUT-X292-LSmitll_DFFT-INt 0 X290-LSmitll_SPLITT-OUT-X292-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X290 X283-LSmitll_NDROT-OUT-X290-LSmitll_SPLITT-IN X290-LSmitll_SPLITT-OUT-X294-LSmitll_NOTT-INt X290-LSmitll_SPLITT-OUT-X292-LSmitll_DFFT-INt LSmitll_SPLITT

t1148 X291-LSmitll_DFFT-OUT-X244-LSmitll_SPLITT-INt 0 X291-LSmitll_DFFT-OUT-X244-LSmitll_SPLITT-IN 0 z0=5 td=3.6ps
X291 X289-LSmitll_SPLITT-OUT-X291-LSmitll_DFFT-IN X511-LSmitll_SPLITT-OUT-X291-LSmitll_DFFT-IN X291-LSmitll_DFFT-OUT-X244-LSmitll_SPLITT-INt LSmitll_DFFT

t1149 X292-LSmitll_DFFT-OUT-X252-LSmitll_XORT-INt 0 X292-LSmitll_DFFT-OUT-X252-LSmitll_XORT-IN 0 z0=5 td=2.9ps
X292 X290-LSmitll_SPLITT-OUT-X292-LSmitll_DFFT-IN X563-LSmitll_SPLITT-OUT-X292-LSmitll_DFFT-IN X292-LSmitll_DFFT-OUT-X252-LSmitll_XORT-INt LSmitll_DFFT

t1150 X293-LSmitll_NOTT-OUT-X296-LSmitll_SPLITT-INt 0 X293-LSmitll_NOTT-OUT-X296-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
X293 X289-LSmitll_SPLITT-OUT-X293-LSmitll_NOTT-IN X564-LSmitll_SPLITT-OUT-X293-LSmitll_NOTT-IN X293-LSmitll_NOTT-OUT-X296-LSmitll_SPLITT-INt LSmitll_NOTT

t1151 X294-LSmitll_NOTT-OUT-X295-LSmitll_SPLITT-INt 0 X294-LSmitll_NOTT-OUT-X295-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X294 X290-LSmitll_SPLITT-OUT-X294-LSmitll_NOTT-IN X565-LSmitll_SPLITT-OUT-X294-LSmitll_NOTT-IN X294-LSmitll_NOTT-OUT-X295-LSmitll_SPLITT-INt LSmitll_NOTT

t1152 X295-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-INt 0 X295-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-IN 0 z0=5 td=3.0ps
t1153 X295-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-INt 0 X295-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-IN 0 z0=5 td=5.8ps
X295 X294-LSmitll_NOTT-OUT-X295-LSmitll_SPLITT-IN X295-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-INt X295-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-INt LSmitll_SPLITT

t1154 X296-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-INt 0 X296-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-IN 0 z0=5 td=5.5ps
t1155 X296-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-INt 0 X296-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-IN 0 z0=5 td=6.5ps
X296 X293-LSmitll_NOTT-OUT-X296-LSmitll_SPLITT-IN X296-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-INt X296-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-INt LSmitll_SPLITT

t1156 X297-LSmitll_DFFT-OUT-X302-LSmitll_DFFT-INt 0 X297-LSmitll_DFFT-OUT-X302-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X297 X285-LSmitll_DFFT-OUT-X297-LSmitll_DFFT-IN X536-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-IN X297-LSmitll_DFFT-OUT-X302-LSmitll_DFFT-INt LSmitll_DFFT

t1157 X298-LSmitll_DFFT-OUT-X301-LSmitll_SPLITT-INt 0 X298-LSmitll_DFFT-OUT-X301-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X298 X286-LSmitll_DFFT-OUT-X298-LSmitll_DFFT-IN X523-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-IN X298-LSmitll_DFFT-OUT-X301-LSmitll_SPLITT-INt LSmitll_DFFT

t1158 X299-LSmitll_DFFT-OUT-X305-LSmitll_DFFT-INt 0 X299-LSmitll_DFFT-OUT-X305-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X299 X287-LSmitll_DFFT-OUT-X299-LSmitll_DFFT-IN X462-LSmitll_SPLITT-OUT-X299-LSmitll_DFFT-IN X299-LSmitll_DFFT-OUT-X305-LSmitll_DFFT-INt LSmitll_DFFT

t1159 X300-LSmitll_DFFT-OUT-X306-LSmitll_DFFT-INt 0 X300-LSmitll_DFFT-OUT-X306-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X300 X288-LSmitll_DFFT-OUT-X300-LSmitll_DFFT-IN X479-LSmitll_SPLITT-OUT-X300-LSmitll_DFFT-IN X300-LSmitll_DFFT-OUT-X306-LSmitll_DFFT-INt LSmitll_DFFT

t1160 X301-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-INt 0 X301-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t1161 X301-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-INt 0 X301-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-IN 0 z0=5 td=3.5ps
X301 X298-LSmitll_DFFT-OUT-X301-LSmitll_SPLITT-IN X301-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-INt X301-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-INt LSmitll_SPLITT


X302 X297-LSmitll_DFFT-OUT-X302-LSmitll_DFFT-IN X537-LSmitll_SPLITT-OUT-X302-LSmitll_DFFT-IN write_flagst LSmitll_DFFT


X303 X301-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-IN X524-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-IN select1t LSmitll_DFFT


X304 X301-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-IN X524-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-IN select0t LSmitll_DFFT

t1165 X305-LSmitll_DFFT-OUT-X307-LSmitll_DFFT-INt 0 X305-LSmitll_DFFT-OUT-X307-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X305 X299-LSmitll_DFFT-OUT-X305-LSmitll_DFFT-IN X462-LSmitll_SPLITT-OUT-X305-LSmitll_DFFT-IN X305-LSmitll_DFFT-OUT-X307-LSmitll_DFFT-INt LSmitll_DFFT

t1166 X306-LSmitll_DFFT-OUT-X308-LSmitll_DFFT-INt 0 X306-LSmitll_DFFT-OUT-X308-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X306 X300-LSmitll_DFFT-OUT-X306-LSmitll_DFFT-IN X469-LSmitll_SPLITT-OUT-X306-LSmitll_DFFT-IN X306-LSmitll_DFFT-OUT-X308-LSmitll_DFFT-INt LSmitll_DFFT

t1167 X307-LSmitll_DFFT-OUT-X309-LSmitll_DFFT-INt 0 X307-LSmitll_DFFT-OUT-X309-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X307 X305-LSmitll_DFFT-OUT-X307-LSmitll_DFFT-IN X463-LSmitll_SPLITT-OUT-X307-LSmitll_DFFT-IN X307-LSmitll_DFFT-OUT-X309-LSmitll_DFFT-INt LSmitll_DFFT

t1168 X308-LSmitll_DFFT-OUT-X310-LSmitll_DFFT-INt 0 X308-LSmitll_DFFT-OUT-X310-LSmitll_DFFT-IN 0 z0=5 td=2.9ps
X308 X306-LSmitll_DFFT-OUT-X308-LSmitll_DFFT-IN X566-LSmitll_SPLITT-OUT-X308-LSmitll_DFFT-IN X308-LSmitll_DFFT-OUT-X310-LSmitll_DFFT-INt LSmitll_DFFT

t1169 X309-LSmitll_DFFT-OUT-X311-LSmitll_OR2T-INt 0 X309-LSmitll_DFFT-OUT-X311-LSmitll_OR2T-IN 0 z0=5 td=2.5ps
X309 X307-LSmitll_DFFT-OUT-X309-LSmitll_DFFT-IN X466-LSmitll_SPLITT-OUT-X309-LSmitll_DFFT-IN X309-LSmitll_DFFT-OUT-X311-LSmitll_OR2T-INt LSmitll_DFFT

t1170 X310-LSmitll_DFFT-OUT-X312-LSmitll_OR2T-INt 0 X310-LSmitll_DFFT-OUT-X312-LSmitll_OR2T-IN 0 z0=5 td=2.5ps
X310 X308-LSmitll_DFFT-OUT-X310-LSmitll_DFFT-IN X480-LSmitll_SPLITT-OUT-X310-LSmitll_DFFT-IN X310-LSmitll_DFFT-OUT-X312-LSmitll_OR2T-INt LSmitll_DFFT


X311 X167-LSmitll_DFFT-OUT-X311-LSmitll_OR2T-IN X309-LSmitll_DFFT-OUT-X311-LSmitll_OR2T-IN X469-LSmitll_SPLITT-OUT-X311-LSmitll_OR2T-IN Addr0t LSmitll_OR2T


X312 X169-LSmitll_DFFT-OUT-X312-LSmitll_OR2T-IN X310-LSmitll_DFFT-OUT-X312-LSmitll_OR2T-IN X480-LSmitll_SPLITT-OUT-X312-LSmitll_OR2T-IN Addr1t LSmitll_OR2T

t1173 X313-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-INt 0 X313-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1174 X313-LSmitll_SPLITT-OUT-X137-LSmitll_AND2T-INt 0 X313-LSmitll_SPLITT-OUT-X137-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
X313 X315-LSmitll_SPLITT-OUT-X313-LSmitll_SPLITT-IN X313-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-INt X313-LSmitll_SPLITT-OUT-X137-LSmitll_AND2T-INt LSmitll_SPLITT

t1175 X314-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-INt 0 X314-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-IN 0 z0=5 td=2.8ps
t1176 X314-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-INt 0 X314-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-IN 0 z0=5 td=3.4ps
X314 X315-LSmitll_SPLITT-OUT-X314-LSmitll_SPLITT-IN X314-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-INt X314-LSmitll_SPLITT-OUT-X93-LSmitll_OR2T-INt LSmitll_SPLITT

t1177 X315-LSmitll_SPLITT-OUT-X313-LSmitll_SPLITT-INt 0 X315-LSmitll_SPLITT-OUT-X313-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
t1178 X315-LSmitll_SPLITT-OUT-X314-LSmitll_SPLITT-INt 0 X315-LSmitll_SPLITT-OUT-X314-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X315 X319-LSmitll_SPLITT-OUT-X315-LSmitll_SPLITT-IN X315-LSmitll_SPLITT-OUT-X313-LSmitll_SPLITT-INt X315-LSmitll_SPLITT-OUT-X314-LSmitll_SPLITT-INt LSmitll_SPLITT

t1179 X316-LSmitll_SPLITT-OUT-X80-LSmitll_NOTT-INt 0 X316-LSmitll_SPLITT-OUT-X80-LSmitll_NOTT-IN 0 z0=5 td=5.9ps
t1180 X316-LSmitll_SPLITT-OUT-X199-LSmitll_DFFT-INt 0 X316-LSmitll_SPLITT-OUT-X199-LSmitll_DFFT-IN 0 z0=5 td=6.3ps
X316 X318-LSmitll_SPLITT-OUT-X316-LSmitll_SPLITT-IN X316-LSmitll_SPLITT-OUT-X80-LSmitll_NOTT-INt X316-LSmitll_SPLITT-OUT-X199-LSmitll_DFFT-INt LSmitll_SPLITT

t1181 X317-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-INt 0 X317-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t1182 X317-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-INt 0 X317-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X317 X318-LSmitll_SPLITT-OUT-X317-LSmitll_SPLITT-IN X317-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-INt X317-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-INt LSmitll_SPLITT

t1183 X318-LSmitll_SPLITT-OUT-X316-LSmitll_SPLITT-INt 0 X318-LSmitll_SPLITT-OUT-X316-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1184 X318-LSmitll_SPLITT-OUT-X317-LSmitll_SPLITT-INt 0 X318-LSmitll_SPLITT-OUT-X317-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X318 X319-LSmitll_SPLITT-OUT-X318-LSmitll_SPLITT-IN X318-LSmitll_SPLITT-OUT-X316-LSmitll_SPLITT-INt X318-LSmitll_SPLITT-OUT-X317-LSmitll_SPLITT-INt LSmitll_SPLITT

t1185 X319-LSmitll_SPLITT-OUT-X315-LSmitll_SPLITT-INt 0 X319-LSmitll_SPLITT-OUT-X315-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1186 X319-LSmitll_SPLITT-OUT-X318-LSmitll_SPLITT-INt 0 X319-LSmitll_SPLITT-OUT-X318-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X319 X326-LSmitll_SPLITT-OUT-X319-LSmitll_SPLITT-IN X319-LSmitll_SPLITT-OUT-X315-LSmitll_SPLITT-INt X319-LSmitll_SPLITT-OUT-X318-LSmitll_SPLITT-INt LSmitll_SPLITT

t1187 X320-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-INt 0 X320-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
t1188 X320-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-INt 0 X320-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
X320 X322-LSmitll_SPLITT-OUT-X320-LSmitll_SPLITT-IN X320-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-INt X320-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-INt LSmitll_SPLITT

t1189 X321-LSmitll_SPLITT-OUT-X141-LSmitll_AND2T-INt 0 X321-LSmitll_SPLITT-OUT-X141-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
t1190 X321-LSmitll_SPLITT-OUT-X157-LSmitll_OR2T-INt 0 X321-LSmitll_SPLITT-OUT-X157-LSmitll_OR2T-IN 0 z0=5 td=1.2ps
X321 X322-LSmitll_SPLITT-OUT-X321-LSmitll_SPLITT-IN X321-LSmitll_SPLITT-OUT-X141-LSmitll_AND2T-INt X321-LSmitll_SPLITT-OUT-X157-LSmitll_OR2T-INt LSmitll_SPLITT

t1191 X322-LSmitll_SPLITT-OUT-X320-LSmitll_SPLITT-INt 0 X322-LSmitll_SPLITT-OUT-X320-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1192 X322-LSmitll_SPLITT-OUT-X321-LSmitll_SPLITT-INt 0 X322-LSmitll_SPLITT-OUT-X321-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X322 X325-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-IN X322-LSmitll_SPLITT-OUT-X320-LSmitll_SPLITT-INt X322-LSmitll_SPLITT-OUT-X321-LSmitll_SPLITT-INt LSmitll_SPLITT

t1193 X323-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-INt 0 X323-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1194 X323-LSmitll_SPLITT-OUT-X224-LSmitll_DFFT-INt 0 X323-LSmitll_SPLITT-OUT-X224-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X323 X324-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-IN X323-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-INt X323-LSmitll_SPLITT-OUT-X224-LSmitll_DFFT-INt LSmitll_SPLITT

t1195 X324-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-INt 0 X324-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1196 X324-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-INt 0 X324-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-IN 0 z0=5 td=1.0ps
X324 X325-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-IN X324-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-INt X324-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-INt LSmitll_SPLITT

t1197 X325-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-INt 0 X325-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1198 X325-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-INt 0 X325-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X325 X326-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-IN X325-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-INt X325-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-INt LSmitll_SPLITT

t1199 X326-LSmitll_SPLITT-OUT-X319-LSmitll_SPLITT-INt 0 X326-LSmitll_SPLITT-OUT-X319-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1200 X326-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-INt 0 X326-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X326 X341-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-IN X326-LSmitll_SPLITT-OUT-X319-LSmitll_SPLITT-INt X326-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-INt LSmitll_SPLITT

t1201 X327-LSmitll_SPLITT-OUT-X185-LSmitll_DFFT-INt 0 X327-LSmitll_SPLITT-OUT-X185-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1202 X327-LSmitll_SPLITT-OUT-X212-LSmitll_DFFT-INt 0 X327-LSmitll_SPLITT-OUT-X212-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
X327 X329-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-IN X327-LSmitll_SPLITT-OUT-X185-LSmitll_DFFT-INt X327-LSmitll_SPLITT-OUT-X212-LSmitll_DFFT-INt LSmitll_SPLITT

t1203 X328-LSmitll_SPLITT-OUT-X125-LSmitll_AND2T-INt 0 X328-LSmitll_SPLITT-OUT-X125-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1204 X328-LSmitll_SPLITT-OUT-X170-LSmitll_DFFT-INt 0 X328-LSmitll_SPLITT-OUT-X170-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X328 X329-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-IN X328-LSmitll_SPLITT-OUT-X125-LSmitll_AND2T-INt X328-LSmitll_SPLITT-OUT-X170-LSmitll_DFFT-INt LSmitll_SPLITT

t1205 X329-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-INt 0 X329-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1206 X329-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-INt 0 X329-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X329 X333-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-IN X329-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-INt X329-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-INt LSmitll_SPLITT

t1207 X330-LSmitll_SPLITT-OUT-X75-LSmitll_DFFT-INt 0 X330-LSmitll_SPLITT-OUT-X75-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
t1208 X330-LSmitll_SPLITT-OUT-X152-LSmitll_OR2T-INt 0 X330-LSmitll_SPLITT-OUT-X152-LSmitll_OR2T-IN 0 z0=5 td=2.1ps
X330 X332-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-IN X330-LSmitll_SPLITT-OUT-X75-LSmitll_DFFT-INt X330-LSmitll_SPLITT-OUT-X152-LSmitll_OR2T-INt LSmitll_SPLITT

t1209 X331-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt 0 X331-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN 0 z0=5 td=1.5ps
t1210 X331-LSmitll_SPLITT-OUT-X153-LSmitll_OR2T-INt 0 X331-LSmitll_SPLITT-OUT-X153-LSmitll_OR2T-IN 0 z0=5 td=3.3ps
X331 X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-IN X331-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt X331-LSmitll_SPLITT-OUT-X153-LSmitll_OR2T-INt LSmitll_SPLITT

t1211 X332-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-INt 0 X332-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1212 X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-INt 0 X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X332 X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-IN X332-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-INt X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-INt LSmitll_SPLITT

t1213 X333-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-INt 0 X333-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-IN 0 z0=5 td=0.5ps
t1214 X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-INt 0 X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X333 X340-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-IN X333-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-INt X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-INt LSmitll_SPLITT

t1215 X334-LSmitll_SPLITT-OUT-X73-LSmitll_DFFT-INt 0 X334-LSmitll_SPLITT-OUT-X73-LSmitll_DFFT-IN 0 z0=5 td=3.9ps
t1216 X334-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-INt 0 X334-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-IN 0 z0=5 td=1.4ps
X334 X336-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-IN X334-LSmitll_SPLITT-OUT-X73-LSmitll_DFFT-INt X334-LSmitll_SPLITT-OUT-X123-LSmitll_AND2T-INt LSmitll_SPLITT

t1217 X335-LSmitll_SPLITT-OUT-X74-LSmitll_DFFT-INt 0 X335-LSmitll_SPLITT-OUT-X74-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
t1218 X335-LSmitll_SPLITT-OUT-X148-LSmitll_DFFT-INt 0 X335-LSmitll_SPLITT-OUT-X148-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
X335 X336-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-IN X335-LSmitll_SPLITT-OUT-X74-LSmitll_DFFT-INt X335-LSmitll_SPLITT-OUT-X148-LSmitll_DFFT-INt LSmitll_SPLITT

t1219 X336-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-INt 0 X336-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1220 X336-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-INt 0 X336-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X336 X339-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-IN X336-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-INt X336-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-INt LSmitll_SPLITT

t1221 X337-LSmitll_SPLITT-OUT-X71-LSmitll_DFFT-INt 0 X337-LSmitll_SPLITT-OUT-X71-LSmitll_DFFT-IN 0 z0=5 td=4.4ps
t1222 X337-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-INt 0 X337-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
X337 X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-IN X337-LSmitll_SPLITT-OUT-X71-LSmitll_DFFT-INt X337-LSmitll_SPLITT-OUT-X127-LSmitll_AND2T-INt LSmitll_SPLITT

t1223 X338-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-INt 0 X338-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1224 X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-INt 0 X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X338 X339-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-IN X338-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-INt X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-INt LSmitll_SPLITT

t1225 X339-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-INt 0 X339-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1226 X339-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-INt 0 X339-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X339 X340-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-IN X339-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-INt X339-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-INt LSmitll_SPLITT

t1227 X340-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-INt 0 X340-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1228 X340-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-INt 0 X340-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-IN 0 z0=5 td=7.5ps
X340 X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-IN X340-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-INt X340-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-INt LSmitll_SPLITT

t1229 X341-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-INt 0 X341-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-IN 0 z0=5 td=6.3ps
t1230 X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-INt 0 X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X341 X370-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-IN X341-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-INt X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-INt LSmitll_SPLITT

t1231 X342-LSmitll_SPLITT-OUT-X140-LSmitll_AND2T-INt 0 X342-LSmitll_SPLITT-OUT-X140-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t1232 X342-LSmitll_SPLITT-OUT-X159-LSmitll_OR2T-INt 0 X342-LSmitll_SPLITT-OUT-X159-LSmitll_OR2T-IN 0 z0=5 td=2.0ps
X342 X344-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-IN X342-LSmitll_SPLITT-OUT-X140-LSmitll_AND2T-INt X342-LSmitll_SPLITT-OUT-X159-LSmitll_OR2T-INt LSmitll_SPLITT

t1233 X343-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-INt 0 X343-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
t1234 X343-LSmitll_SPLITT-OUT-X139-LSmitll_AND2T-INt 0 X343-LSmitll_SPLITT-OUT-X139-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
X343 X344-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-IN X343-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-INt X343-LSmitll_SPLITT-OUT-X139-LSmitll_AND2T-INt LSmitll_SPLITT

t1235 X344-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-INt 0 X344-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1236 X344-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-INt 0 X344-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X344 X348-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-IN X344-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-INt X344-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-INt LSmitll_SPLITT

t1237 X345-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-INt 0 X345-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-IN 0 z0=5 td=2.8ps
t1238 X345-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-INt 0 X345-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
X345 X347-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-IN X345-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-INt X345-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-INt LSmitll_SPLITT

t1239 X346-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-INt 0 X346-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
t1240 X346-LSmitll_SPLITT-OUT-X192-LSmitll_OR2T-INt 0 X346-LSmitll_SPLITT-OUT-X192-LSmitll_OR2T-IN 0 z0=5 td=2.0ps
X346 X347-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-IN X346-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-INt X346-LSmitll_SPLITT-OUT-X192-LSmitll_OR2T-INt LSmitll_SPLITT

t1241 X347-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-INt 0 X347-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-IN 0 z0=5 td=1.0ps
t1242 X347-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-INt 0 X347-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X347 X348-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-IN X347-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-INt X347-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-INt LSmitll_SPLITT

t1243 X348-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-INt 0 X348-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
t1244 X348-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-INt 0 X348-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X348 X355-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-IN X348-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-INt X348-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-INt LSmitll_SPLITT

t1245 X349-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-INt 0 X349-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
t1246 X349-LSmitll_SPLITT-OUT-X158-LSmitll_OR2T-INt 0 X349-LSmitll_SPLITT-OUT-X158-LSmitll_OR2T-IN 0 z0=5 td=0.8ps
X349 X351-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-IN X349-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-INt X349-LSmitll_SPLITT-OUT-X158-LSmitll_OR2T-INt LSmitll_SPLITT

t1247 X350-LSmitll_SPLITT-OUT-X35-LSmitll_XORT-INt 0 X350-LSmitll_SPLITT-OUT-X35-LSmitll_XORT-IN 0 z0=5 td=2.1ps
t1248 X350-LSmitll_SPLITT-OUT-X90-LSmitll_AND2T-INt 0 X350-LSmitll_SPLITT-OUT-X90-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X350 X351-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-IN X350-LSmitll_SPLITT-OUT-X35-LSmitll_XORT-INt X350-LSmitll_SPLITT-OUT-X90-LSmitll_AND2T-INt LSmitll_SPLITT

t1249 X351-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-INt 0 X351-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1250 X351-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-INt 0 X351-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X351 X354-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-IN X351-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-INt X351-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-INt LSmitll_SPLITT

t1251 X352-LSmitll_SPLITT-OUT-X149-LSmitll_DFFT-INt 0 X352-LSmitll_SPLITT-OUT-X149-LSmitll_DFFT-IN 0 z0=5 td=3.3ps
t1252 X352-LSmitll_SPLITT-OUT-X176-LSmitll_OR2T-INt 0 X352-LSmitll_SPLITT-OUT-X176-LSmitll_OR2T-IN 0 z0=5 td=0.6ps
X352 X353-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-IN X352-LSmitll_SPLITT-OUT-X149-LSmitll_DFFT-INt X352-LSmitll_SPLITT-OUT-X176-LSmitll_OR2T-INt LSmitll_SPLITT

t1253 X353-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-INt 0 X353-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1254 X353-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-INt 0 X353-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X353 X354-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-IN X353-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-INt X353-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-INt LSmitll_SPLITT

t1255 X354-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-INt 0 X354-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
t1256 X354-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-INt 0 X354-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X354 X355-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-IN X354-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-INt X354-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-INt LSmitll_SPLITT

t1257 X355-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-INt 0 X355-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1258 X355-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-INt 0 X355-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X355 X369-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-IN X355-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-INt X355-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-INt LSmitll_SPLITT

t1259 X356-LSmitll_SPLITT-OUT-X248-LSmitll_DFFT-INt 0 X356-LSmitll_SPLITT-OUT-X248-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
t1260 X356-LSmitll_SPLITT-OUT-X256-LSmitll_DFFT-INt 0 X356-LSmitll_SPLITT-OUT-X256-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
X356 X358-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-IN X356-LSmitll_SPLITT-OUT-X248-LSmitll_DFFT-INt X356-LSmitll_SPLITT-OUT-X256-LSmitll_DFFT-INt LSmitll_SPLITT

t1261 X357-LSmitll_SPLITT-OUT-X69-LSmitll_NOTT-INt 0 X357-LSmitll_SPLITT-OUT-X69-LSmitll_NOTT-IN 0 z0=5 td=1.0ps
t1262 X357-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt 0 X357-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
X357 X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-IN X357-LSmitll_SPLITT-OUT-X69-LSmitll_NOTT-INt X357-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt LSmitll_SPLITT

t1263 X358-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-INt 0 X358-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1264 X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-INt 0 X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X358 X361-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-IN X358-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-INt X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-INt LSmitll_SPLITT

t1265 X359-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-INt 0 X359-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
t1266 X359-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-INt 0 X359-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X359 X360-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-IN X359-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-INt X359-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-INt LSmitll_SPLITT

t1267 X360-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-INt 0 X360-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1268 X360-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-INt 0 X360-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X360 X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-IN X360-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-INt X360-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-INt LSmitll_SPLITT

t1269 X361-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-INt 0 X361-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1270 X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-INt 0 X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-IN 0 z0=5 td=4.2ps
X361 X368-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-IN X361-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-INt X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-INt LSmitll_SPLITT

t1271 X362-LSmitll_SPLITT-OUT-X70-LSmitll_DFFT-INt 0 X362-LSmitll_SPLITT-OUT-X70-LSmitll_DFFT-IN 0 z0=5 td=3.9ps
t1272 X362-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-INt 0 X362-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
X362 X364-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-IN X362-LSmitll_SPLITT-OUT-X70-LSmitll_DFFT-INt X362-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-INt LSmitll_SPLITT

t1273 X363-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-INt 0 X363-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-IN 0 z0=5 td=0.7ps
t1274 X363-LSmitll_SPLITT-OUT-X213-LSmitll_DFFT-INt 0 X363-LSmitll_SPLITT-OUT-X213-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
X363 X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-IN X363-LSmitll_SPLITT-OUT-X119-LSmitll_AND2T-INt X363-LSmitll_SPLITT-OUT-X213-LSmitll_DFFT-INt LSmitll_SPLITT

t1275 X364-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-INt 0 X364-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1276 X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-INt 0 X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X364 X367-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-IN X364-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-INt X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-INt LSmitll_SPLITT

t1277 X365-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-INt 0 X365-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-IN 0 z0=5 td=2.5ps
t1278 X365-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-INt 0 X365-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-IN 0 z0=5 td=2.9ps
X365 X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-IN X365-LSmitll_SPLITT-OUT-X117-LSmitll_OR2T-INt X365-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-INt LSmitll_SPLITT

t1279 X366-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-INt 0 X366-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1280 X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-INt 0 X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X366 X367-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-IN X366-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-INt X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-INt LSmitll_SPLITT

t1281 X367-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-INt 0 X367-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1282 X367-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-INt 0 X367-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X367 X368-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-IN X367-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-INt X367-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-INt LSmitll_SPLITT

t1283 X368-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-INt 0 X368-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
t1284 X368-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-INt 0 X368-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X368 X369-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-IN X368-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-INt X368-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-INt LSmitll_SPLITT

t1285 X369-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-INt 0 X369-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-IN 0 z0=5 td=4.3ps
t1286 X369-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-INt 0 X369-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X369 X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-IN X369-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-INt X369-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-INt LSmitll_SPLITT

t1287 X370-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-INt 0 X370-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-IN 0 z0=5 td=5.7ps
t1288 X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-INt 0 X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-IN 0 z0=5 td=5.2ps
X370 X429-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-IN X370-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-INt X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-INt LSmitll_SPLITT

t1289 X371-LSmitll_SPLITT-OUT-X171-LSmitll_DFFT-INt 0 X371-LSmitll_SPLITT-OUT-X171-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t1290 X371-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-INt 0 X371-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-IN 0 z0=5 td=0.3ps
X371 X373-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-IN X371-LSmitll_SPLITT-OUT-X171-LSmitll_DFFT-INt X371-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-INt LSmitll_SPLITT

t1291 X372-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-INt 0 X372-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1292 X372-LSmitll_SPLITT-OUT-X179-LSmitll_DFFT-INt 0 X372-LSmitll_SPLITT-OUT-X179-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
X372 X373-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-IN X372-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-INt X372-LSmitll_SPLITT-OUT-X179-LSmitll_DFFT-INt LSmitll_SPLITT

t1293 X373-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-INt 0 X373-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1294 X373-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-INt 0 X373-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X373 X377-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-IN X373-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-INt X373-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-INt LSmitll_SPLITT

t1295 X374-LSmitll_SPLITT-OUT-X194-LSmitll_DFFT-INt 0 X374-LSmitll_SPLITT-OUT-X194-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
t1296 X374-LSmitll_SPLITT-OUT-X205-LSmitll_DFFT-INt 0 X374-LSmitll_SPLITT-OUT-X205-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
X374 X376-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-IN X374-LSmitll_SPLITT-OUT-X194-LSmitll_DFFT-INt X374-LSmitll_SPLITT-OUT-X205-LSmitll_DFFT-INt LSmitll_SPLITT

t1297 X375-LSmitll_SPLITT-OUT-X219-LSmitll_AND2T-INt 0 X375-LSmitll_SPLITT-OUT-X219-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
t1298 X375-LSmitll_SPLITT-OUT-X233-LSmitll_OR2T-INt 0 X375-LSmitll_SPLITT-OUT-X233-LSmitll_OR2T-IN 0 z0=5 td=0.9ps
X375 X376-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-IN X375-LSmitll_SPLITT-OUT-X219-LSmitll_AND2T-INt X375-LSmitll_SPLITT-OUT-X233-LSmitll_OR2T-INt LSmitll_SPLITT

t1299 X376-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-INt 0 X376-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1300 X376-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-INt 0 X376-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X376 X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-IN X376-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-INt X376-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-INt LSmitll_SPLITT

t1301 X377-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-INt 0 X377-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1302 X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-INt 0 X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X377 X384-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-IN X377-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-INt X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-INt LSmitll_SPLITT

t1303 X378-LSmitll_SPLITT-OUT-X135-LSmitll_OR2T-INt 0 X378-LSmitll_SPLITT-OUT-X135-LSmitll_OR2T-IN 0 z0=5 td=2.1ps
t1304 X378-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-INt 0 X378-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
X378 X380-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-IN X378-LSmitll_SPLITT-OUT-X135-LSmitll_OR2T-INt X378-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-INt LSmitll_SPLITT

t1305 X379-LSmitll_SPLITT-OUT-X76-LSmitll_DFFT-INt 0 X379-LSmitll_SPLITT-OUT-X76-LSmitll_DFFT-IN 0 z0=5 td=2.8ps
t1306 X379-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-INt 0 X379-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
X379 X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-IN X379-LSmitll_SPLITT-OUT-X76-LSmitll_DFFT-INt X379-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-INt LSmitll_SPLITT

t1307 X380-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-INt 0 X380-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1308 X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-INt 0 X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X380 X383-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-IN X380-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-INt X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-INt LSmitll_SPLITT

t1309 X381-LSmitll_SPLITT-OUT-X191-LSmitll_DFFT-INt 0 X381-LSmitll_SPLITT-OUT-X191-LSmitll_DFFT-IN 0 z0=5 td=2.8ps
t1310 X381-LSmitll_SPLITT-OUT-X220-LSmitll_DFFT-INt 0 X381-LSmitll_SPLITT-OUT-X220-LSmitll_DFFT-IN 0 z0=5 td=4.5ps
X381 X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-IN X381-LSmitll_SPLITT-OUT-X191-LSmitll_DFFT-INt X381-LSmitll_SPLITT-OUT-X220-LSmitll_DFFT-INt LSmitll_SPLITT

t1311 X382-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-INt 0 X382-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-IN 0 z0=5 td=3.4ps
t1312 X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-INt 0 X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X382 X383-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-IN X382-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-INt X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-INt LSmitll_SPLITT

t1313 X383-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-INt 0 X383-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t1314 X383-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-INt 0 X383-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X383 X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-IN X383-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-INt X383-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-INt LSmitll_SPLITT

t1315 X384-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-INt 0 X384-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1316 X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-INt 0 X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X384 X399-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-IN X384-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-INt X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-INt LSmitll_SPLITT

t1317 X385-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-INt 0 X385-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1318 X385-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-INt 0 X385-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-IN 0 z0=5 td=3.0ps
X385 X387-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-IN X385-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-INt X385-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-INt LSmitll_SPLITT

t1319 X386-LSmitll_SPLITT-OUT-X215-LSmitll_DFFT-INt 0 X386-LSmitll_SPLITT-OUT-X215-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
t1320 X386-LSmitll_SPLITT-OUT-X227-LSmitll_DFFT-INt 0 X386-LSmitll_SPLITT-OUT-X227-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
X386 X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-IN X386-LSmitll_SPLITT-OUT-X215-LSmitll_DFFT-INt X386-LSmitll_SPLITT-OUT-X227-LSmitll_DFFT-INt LSmitll_SPLITT

t1321 X387-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-INt 0 X387-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-IN 0 z0=5 td=1.0ps
t1322 X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-INt 0 X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
X387 X391-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-IN X387-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-INt X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-INt LSmitll_SPLITT

t1323 X388-LSmitll_SPLITT-OUT-X231-LSmitll_DFFT-INt 0 X388-LSmitll_SPLITT-OUT-X231-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t1324 X388-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-INt 0 X388-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
X388 X390-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-IN X388-LSmitll_SPLITT-OUT-X231-LSmitll_DFFT-INt X388-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-INt LSmitll_SPLITT

t1325 X389-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-INt 0 X389-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
t1326 X389-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-INt 0 X389-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-IN 0 z0=5 td=3.3ps
X389 X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-IN X389-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-INt X389-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-INt LSmitll_SPLITT

t1327 X390-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-INt 0 X390-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1328 X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-INt 0 X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X390 X391-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-IN X390-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-INt X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-INt LSmitll_SPLITT

t1329 X391-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-INt 0 X391-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-IN 0 z0=5 td=3.5ps
t1330 X391-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-INt 0 X391-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X391 X398-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-IN X391-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-INt X391-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-INt LSmitll_SPLITT

t1331 X392-LSmitll_SPLITT-OUT-X253-LSmitll_OR2T-INt 0 X392-LSmitll_SPLITT-OUT-X253-LSmitll_OR2T-IN 0 z0=5 td=2.5ps
t1332 X392-LSmitll_SPLITT-OUT-X283-LSmitll_NDROT-INt 0 X392-LSmitll_SPLITT-OUT-X283-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
X392 X394-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-IN X392-LSmitll_SPLITT-OUT-X253-LSmitll_OR2T-INt X392-LSmitll_SPLITT-OUT-X283-LSmitll_NDROT-INt LSmitll_SPLITT

t1333 X393-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-INt 0 X393-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
t1334 X393-LSmitll_SPLITT-OUT-X240-LSmitll_OR2T-INt 0 X393-LSmitll_SPLITT-OUT-X240-LSmitll_OR2T-IN 0 z0=5 td=2.4ps
X393 X394-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-IN X393-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-INt X393-LSmitll_SPLITT-OUT-X240-LSmitll_OR2T-INt LSmitll_SPLITT

t1335 X394-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-INt 0 X394-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1336 X394-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-INt 0 X394-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X394 X397-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-IN X394-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-INt X394-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-INt LSmitll_SPLITT

t1337 X395-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-INt 0 X395-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-IN 0 z0=5 td=0.4ps
t1338 X395-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-INt 0 X395-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-IN 0 z0=5 td=1.5ps
X395 X396-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-IN X395-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-INt X395-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-INt LSmitll_SPLITT

t1339 X396-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-INt 0 X396-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-IN 0 z0=5 td=1.0ps
t1340 X396-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-INt 0 X396-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X396 X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-IN X396-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-INt X396-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-INt LSmitll_SPLITT

t1341 X397-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-INt 0 X397-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1342 X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-INt 0 X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X397 X398-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-IN X397-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-INt X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-INt LSmitll_SPLITT

t1343 X398-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-INt 0 X398-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1344 X398-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-INt 0 X398-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
X398 X399-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-IN X398-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-INt X398-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-INt LSmitll_SPLITT

t1345 X399-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-INt 0 X399-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
t1346 X399-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-INt 0 X399-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X399 X428-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-IN X399-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-INt X399-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-INt LSmitll_SPLITT

t1347 X400-LSmitll_SPLITT-OUT-X72-LSmitll_DFFT-INt 0 X400-LSmitll_SPLITT-OUT-X72-LSmitll_DFFT-IN 0 z0=5 td=0.4ps
t1348 X400-LSmitll_SPLITT-OUT-X115-LSmitll_DFFT-INt 0 X400-LSmitll_SPLITT-OUT-X115-LSmitll_DFFT-IN 0 z0=5 td=1.7ps
X400 X402-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-IN X400-LSmitll_SPLITT-OUT-X72-LSmitll_DFFT-INt X400-LSmitll_SPLITT-OUT-X115-LSmitll_DFFT-INt LSmitll_SPLITT

t1349 X401-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-INt 0 X401-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-IN 0 z0=5 td=3.4ps
t1350 X401-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-INt 0 X401-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-IN 0 z0=5 td=3.4ps
X401 X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-IN X401-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-INt X401-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-INt LSmitll_SPLITT

t1351 X402-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-INt 0 X402-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1352 X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-INt 0 X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
X402 X406-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-IN X402-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-INt X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-INt LSmitll_SPLITT

t1353 X403-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-INt 0 X403-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
t1354 X403-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-INt 0 X403-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-IN 0 z0=5 td=1.9ps
X403 X405-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-IN X403-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-INt X403-LSmitll_SPLITT-OUT-X202-LSmitll_AND2T-INt LSmitll_SPLITT

t1355 X404-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-INt 0 X404-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-IN 0 z0=5 td=4.4ps
t1356 X404-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-INt 0 X404-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-IN 0 z0=5 td=3.1ps
X404 X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-IN X404-LSmitll_SPLITT-OUT-X129-LSmitll_AND2T-INt X404-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-INt LSmitll_SPLITT

t1357 X405-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-INt 0 X405-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1358 X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-INt 0 X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X405 X406-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-IN X405-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-INt X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-INt LSmitll_SPLITT

t1359 X406-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-INt 0 X406-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1360 X406-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-INt 0 X406-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
X406 X413-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-IN X406-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-INt X406-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-INt LSmitll_SPLITT

t1361 X407-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-INt 0 X407-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t1362 X407-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-INt 0 X407-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
X407 X409-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-IN X407-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-INt X407-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-INt LSmitll_SPLITT

t1363 X408-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-INt 0 X408-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1364 X408-LSmitll_SPLITT-OUT-X197-LSmitll_DFFT-INt 0 X408-LSmitll_SPLITT-OUT-X197-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
X408 X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-IN X408-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-INt X408-LSmitll_SPLITT-OUT-X197-LSmitll_DFFT-INt LSmitll_SPLITT

t1365 X409-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-INt 0 X409-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1366 X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-INt 0 X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X409 X412-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-IN X409-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-INt X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-INt LSmitll_SPLITT

t1367 X410-LSmitll_SPLITT-OUT-X203-LSmitll_NOTT-INt 0 X410-LSmitll_SPLITT-OUT-X203-LSmitll_NOTT-IN 0 z0=5 td=1.1ps
t1368 X410-LSmitll_SPLITT-OUT-X214-LSmitll_AND2T-INt 0 X410-LSmitll_SPLITT-OUT-X214-LSmitll_AND2T-IN 0 z0=5 td=1.3ps
X410 X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-IN X410-LSmitll_SPLITT-OUT-X203-LSmitll_NOTT-INt X410-LSmitll_SPLITT-OUT-X214-LSmitll_AND2T-INt LSmitll_SPLITT

t1369 X411-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-INt 0 X411-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-IN 0 z0=5 td=2.8ps
t1370 X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-INt 0 X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-IN 0 z0=5 td=0.6ps
X411 X412-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-IN X411-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-INt X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-INt LSmitll_SPLITT

t1371 X412-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-INt 0 X412-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1372 X412-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-INt 0 X412-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X412 X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-IN X412-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-INt X412-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-INt LSmitll_SPLITT

t1373 X413-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-INt 0 X413-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1374 X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-INt 0 X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-IN 0 z0=5 td=3.4ps
X413 X427-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-IN X413-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-INt X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-INt LSmitll_SPLITT

t1375 X414-LSmitll_SPLITT-OUT-X229-LSmitll_AND2T-INt 0 X414-LSmitll_SPLITT-OUT-X229-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1376 X414-LSmitll_SPLITT-OUT-X252-LSmitll_XORT-INt 0 X414-LSmitll_SPLITT-OUT-X252-LSmitll_XORT-IN 0 z0=5 td=4.2ps
X414 X416-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-IN X414-LSmitll_SPLITT-OUT-X229-LSmitll_AND2T-INt X414-LSmitll_SPLITT-OUT-X252-LSmitll_XORT-INt LSmitll_SPLITT

t1377 X415-LSmitll_SPLITT-OUT-X217-LSmitll_DFFT-INt 0 X415-LSmitll_SPLITT-OUT-X217-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
t1378 X415-LSmitll_SPLITT-OUT-X243-LSmitll_AND2T-INt 0 X415-LSmitll_SPLITT-OUT-X243-LSmitll_AND2T-IN 0 z0=5 td=1.3ps
X415 X416-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-IN X415-LSmitll_SPLITT-OUT-X217-LSmitll_DFFT-INt X415-LSmitll_SPLITT-OUT-X243-LSmitll_AND2T-INt LSmitll_SPLITT

t1379 X416-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-INt 0 X416-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1380 X416-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-INt 0 X416-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
X416 X419-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-IN X416-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-INt X416-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-INt LSmitll_SPLITT

t1381 X417-LSmitll_SPLITT-OUT-X259-LSmitll_XORT-INt 0 X417-LSmitll_SPLITT-OUT-X259-LSmitll_XORT-IN 0 z0=5 td=2.6ps
t1382 X417-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-INt 0 X417-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-IN 0 z0=5 td=2.9ps
X417 X418-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-IN X417-LSmitll_SPLITT-OUT-X259-LSmitll_XORT-INt X417-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-INt LSmitll_SPLITT

t1383 X418-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-INt 0 X418-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-IN 0 z0=5 td=3.7ps
t1384 X418-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-INt 0 X418-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X418 X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-IN X418-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-INt X418-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-INt LSmitll_SPLITT

t1385 X419-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-INt 0 X419-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t1386 X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-INt 0 X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X419 X426-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-IN X419-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-INt X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-INt LSmitll_SPLITT

t1387 X420-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-INt 0 X420-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-IN 0 z0=5 td=1.5ps
t1388 X420-LSmitll_SPLITT-OUT-X230-LSmitll_OR2T-INt 0 X420-LSmitll_SPLITT-OUT-X230-LSmitll_OR2T-IN 0 z0=5 td=1.8ps
X420 X422-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-IN X420-LSmitll_SPLITT-OUT-X216-LSmitll_OR2T-INt X420-LSmitll_SPLITT-OUT-X230-LSmitll_OR2T-INt LSmitll_SPLITT

t1389 X421-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-INt 0 X421-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-IN 0 z0=5 td=1.8ps
t1390 X421-LSmitll_SPLITT-OUT-X241-LSmitll_OR2T-INt 0 X421-LSmitll_SPLITT-OUT-X241-LSmitll_OR2T-IN 0 z0=5 td=0.6ps
X421 X422-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-IN X421-LSmitll_SPLITT-OUT-X232-LSmitll_OR2T-INt X421-LSmitll_SPLITT-OUT-X241-LSmitll_OR2T-INt LSmitll_SPLITT

t1391 X422-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-INt 0 X422-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1392 X422-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-INt 0 X422-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X422 X425-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-IN X422-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-INt X422-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-INt LSmitll_SPLITT

t1393 X423-LSmitll_SPLITT-OUT-X273-LSmitll_DFFT-INt 0 X423-LSmitll_SPLITT-OUT-X273-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
t1394 X423-LSmitll_SPLITT-OUT-X275-LSmitll_DFFT-INt 0 X423-LSmitll_SPLITT-OUT-X275-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X423 X424-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-IN X423-LSmitll_SPLITT-OUT-X273-LSmitll_DFFT-INt X423-LSmitll_SPLITT-OUT-X275-LSmitll_DFFT-INt LSmitll_SPLITT

t1395 X424-LSmitll_SPLITT-OUT-X565-LSmitll_SPLITT-INt 0 X424-LSmitll_SPLITT-OUT-X565-LSmitll_SPLITT-IN 0 z0=5 td=3.2ps
t1396 X424-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-INt 0 X424-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X424 X425-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-IN X424-LSmitll_SPLITT-OUT-X565-LSmitll_SPLITT-INt X424-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-INt LSmitll_SPLITT

t1397 X425-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-INt 0 X425-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1398 X425-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-INt 0 X425-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X425 X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-IN X425-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-INt X425-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-INt LSmitll_SPLITT

t1399 X426-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-INt 0 X426-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
t1400 X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-INt 0 X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X426 X427-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-IN X426-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-INt X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-INt LSmitll_SPLITT

t1401 X427-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-INt 0 X427-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
t1402 X427-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-INt 0 X427-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
X427 X428-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-IN X427-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-INt X427-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-INt LSmitll_SPLITT

t1403 X428-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-INt 0 X428-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
t1404 X428-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-INt 0 X428-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-IN 0 z0=5 td=3.7ps
X428 X429-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-IN X428-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-INt X428-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-INt LSmitll_SPLITT

t1405 X429-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-INt 0 X429-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-IN 0 z0=5 td=5.3ps
t1406 X429-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-INt 0 X429-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-IN 0 z0=5 td=6.8ps
X429 X567-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-IN X429-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-INt X429-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-INt LSmitll_SPLITT

t1407 X430-LSmitll_SPLITT-OUT-X15-LSmitll_DFFT-INt 0 X430-LSmitll_SPLITT-OUT-X15-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1408 X430-LSmitll_SPLITT-OUT-X138-LSmitll_AND2T-INt 0 X430-LSmitll_SPLITT-OUT-X138-LSmitll_AND2T-IN 0 z0=5 td=3.0ps
X430 X432-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-IN X430-LSmitll_SPLITT-OUT-X15-LSmitll_DFFT-INt X430-LSmitll_SPLITT-OUT-X138-LSmitll_AND2T-INt LSmitll_SPLITT

t1409 X431-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-INt 0 X431-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-IN 0 z0=5 td=0.6ps
t1410 X431-LSmitll_SPLITT-OUT-X83-LSmitll_DFFT-INt 0 X431-LSmitll_SPLITT-OUT-X83-LSmitll_DFFT-IN 0 z0=5 td=5.2ps
X431 X432-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-IN X431-LSmitll_SPLITT-OUT-X19-LSmitll_XORT-INt X431-LSmitll_SPLITT-OUT-X83-LSmitll_DFFT-INt LSmitll_SPLITT

t1411 X432-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-INt 0 X432-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1412 X432-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-INt 0 X432-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X432 X436-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-IN X432-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-INt X432-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-INt LSmitll_SPLITT

t1413 X433-LSmitll_SPLITT-OUT-X9-LSmitll_DFFT-INt 0 X433-LSmitll_SPLITT-OUT-X9-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
t1414 X433-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-INt 0 X433-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
X433 X435-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-IN X433-LSmitll_SPLITT-OUT-X9-LSmitll_DFFT-INt X433-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-INt LSmitll_SPLITT

t1415 X434-LSmitll_SPLITT-OUT-X8-LSmitll_DFFT-INt 0 X434-LSmitll_SPLITT-OUT-X8-LSmitll_DFFT-IN 0 z0=5 td=3.2ps
t1416 X434-LSmitll_SPLITT-OUT-X84-LSmitll_NOTT-INt 0 X434-LSmitll_SPLITT-OUT-X84-LSmitll_NOTT-IN 0 z0=5 td=1.8ps
X434 X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-IN X434-LSmitll_SPLITT-OUT-X8-LSmitll_DFFT-INt X434-LSmitll_SPLITT-OUT-X84-LSmitll_NOTT-INt LSmitll_SPLITT

t1417 X435-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-INt 0 X435-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
t1418 X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-INt 0 X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X435 X436-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-IN X435-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-INt X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-INt LSmitll_SPLITT

t1419 X436-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-INt 0 X436-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1420 X436-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-INt 0 X436-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X436 X443-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-IN X436-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-INt X436-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-INt LSmitll_SPLITT

t1421 X437-LSmitll_SPLITT-OUT-X7-LSmitll_DFFT-INt 0 X437-LSmitll_SPLITT-OUT-X7-LSmitll_DFFT-IN 0 z0=5 td=3.2ps
t1422 X437-LSmitll_SPLITT-OUT-X36-LSmitll_NOTT-INt 0 X437-LSmitll_SPLITT-OUT-X36-LSmitll_NOTT-IN 0 z0=5 td=1.9ps
X437 X439-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-IN X437-LSmitll_SPLITT-OUT-X7-LSmitll_DFFT-INt X437-LSmitll_SPLITT-OUT-X36-LSmitll_NOTT-INt LSmitll_SPLITT

t1423 X438-LSmitll_SPLITT-OUT-X16-LSmitll_DFFT-INt 0 X438-LSmitll_SPLITT-OUT-X16-LSmitll_DFFT-IN 0 z0=5 td=1.8ps
t1424 X438-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-INt 0 X438-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X438 X439-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-IN X438-LSmitll_SPLITT-OUT-X16-LSmitll_DFFT-INt X438-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-INt LSmitll_SPLITT

t1425 X439-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-INt 0 X439-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1426 X439-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-INt 0 X439-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X439 X442-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-IN X439-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-INt X439-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-INt LSmitll_SPLITT

t1427 X440-LSmitll_SPLITT-OUT-X249-LSmitll_DFFT-INt 0 X440-LSmitll_SPLITT-OUT-X249-LSmitll_DFFT-IN 0 z0=5 td=3.0ps
t1428 X440-LSmitll_SPLITT-OUT-X271-LSmitll_DFFT-INt 0 X440-LSmitll_SPLITT-OUT-X271-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X440 X441-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-IN X440-LSmitll_SPLITT-OUT-X249-LSmitll_DFFT-INt X440-LSmitll_SPLITT-OUT-X271-LSmitll_DFFT-INt LSmitll_SPLITT

t1429 X441-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-INt 0 X441-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1430 X441-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-INt 0 X441-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X441 X442-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-IN X441-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-INt X441-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-INt LSmitll_SPLITT

t1431 X442-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-INt 0 X442-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1432 X442-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-INt 0 X442-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X442 X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-IN X442-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-INt X442-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-INt LSmitll_SPLITT

t1433 X443-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-INt 0 X443-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
t1434 X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-INt 0 X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X443 X458-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-IN X443-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-INt X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-INt LSmitll_SPLITT

t1435 X444-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-INt 0 X444-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1436 X444-LSmitll_SPLITT-OUT-X200-LSmitll_DFFT-INt 0 X444-LSmitll_SPLITT-OUT-X200-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
X444 X446-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-IN X444-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-INt X444-LSmitll_SPLITT-OUT-X200-LSmitll_DFFT-INt LSmitll_SPLITT

t1437 X445-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-INt 0 X445-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1438 X445-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-INt 0 X445-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X445 X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-IN X445-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-INt X445-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-INt LSmitll_SPLITT

t1439 X446-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-INt 0 X446-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1440 X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-INt 0 X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X446 X450-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-IN X446-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-INt X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-INt LSmitll_SPLITT

t1441 X447-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-INt 0 X447-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-IN 0 z0=5 td=2.8ps
t1442 X447-LSmitll_SPLITT-OUT-X168-LSmitll_DFFT-INt 0 X447-LSmitll_SPLITT-OUT-X168-LSmitll_DFFT-IN 0 z0=5 td=5.8ps
X447 X449-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-IN X447-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-INt X447-LSmitll_SPLITT-OUT-X168-LSmitll_DFFT-INt LSmitll_SPLITT

t1443 X448-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-INt 0 X448-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-IN 0 z0=5 td=3.3ps
t1444 X448-LSmitll_SPLITT-OUT-X150-LSmitll_DFFT-INt 0 X448-LSmitll_SPLITT-OUT-X150-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
X448 X449-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-IN X448-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-INt X448-LSmitll_SPLITT-OUT-X150-LSmitll_DFFT-INt LSmitll_SPLITT

t1445 X449-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-INt 0 X449-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1446 X449-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-INt 0 X449-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
X449 X450-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-IN X449-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-INt X449-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-INt LSmitll_SPLITT

t1447 X450-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-INt 0 X450-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1448 X450-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-INt 0 X450-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X450 X457-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-IN X450-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-INt X450-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-INt LSmitll_SPLITT

t1449 X451-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-INt 0 X451-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1450 X451-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt 0 X451-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN 0 z0=5 td=2.6ps
X451 X453-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-IN X451-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-INt X451-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt LSmitll_SPLITT

t1451 X452-LSmitll_SPLITT-OUT-X3-LSmitll_DFFT-INt 0 X452-LSmitll_SPLITT-OUT-X3-LSmitll_DFFT-IN 0 z0=5 td=2.9ps
t1452 X452-LSmitll_SPLITT-OUT-X257-LSmitll_DFFT-INt 0 X452-LSmitll_SPLITT-OUT-X257-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
X452 X453-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-IN X452-LSmitll_SPLITT-OUT-X3-LSmitll_DFFT-INt X452-LSmitll_SPLITT-OUT-X257-LSmitll_DFFT-INt LSmitll_SPLITT

t1453 X453-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-INt 0 X453-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1454 X453-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-INt 0 X453-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X453 X456-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-IN X453-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-INt X453-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-INt LSmitll_SPLITT

t1455 X454-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-INt 0 X454-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1456 X454-LSmitll_SPLITT-OUT-X118-LSmitll_DFFT-INt 0 X454-LSmitll_SPLITT-OUT-X118-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X454 X455-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-IN X454-LSmitll_SPLITT-OUT-X27-LSmitll_AND2T-INt X454-LSmitll_SPLITT-OUT-X118-LSmitll_DFFT-INt LSmitll_SPLITT

t1457 X455-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-INt 0 X455-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1458 X455-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-INt 0 X455-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X455 X456-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-IN X455-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-INt X455-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-INt LSmitll_SPLITT

t1459 X456-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-INt 0 X456-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1460 X456-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-INt 0 X456-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X456 X457-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-IN X456-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-INt X456-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-INt LSmitll_SPLITT

t1461 X457-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-INt 0 X457-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1462 X457-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-INt 0 X457-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-IN 0 z0=5 td=3.2ps
X457 X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-IN X457-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-INt X457-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-INt LSmitll_SPLITT

t1463 X458-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-INt 0 X458-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-IN 0 z0=5 td=4.0ps
t1464 X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-INt 0 X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
X458 X487-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-IN X458-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-INt X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-INt LSmitll_SPLITT

t1465 X459-LSmitll_SPLITT-OUT-X10-LSmitll_DFFT-INt 0 X459-LSmitll_SPLITT-OUT-X10-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
t1466 X459-LSmitll_SPLITT-OUT-X87-LSmitll_DFFT-INt 0 X459-LSmitll_SPLITT-OUT-X87-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
X459 X461-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-IN X459-LSmitll_SPLITT-OUT-X10-LSmitll_DFFT-INt X459-LSmitll_SPLITT-OUT-X87-LSmitll_DFFT-INt LSmitll_SPLITT

t1467 X460-LSmitll_SPLITT-OUT-X17-LSmitll_NOTT-INt 0 X460-LSmitll_SPLITT-OUT-X17-LSmitll_NOTT-IN 0 z0=5 td=2.0ps
t1468 X460-LSmitll_SPLITT-OUT-X88-LSmitll_NOTT-INt 0 X460-LSmitll_SPLITT-OUT-X88-LSmitll_NOTT-IN 0 z0=5 td=0.9ps
X460 X461-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-IN X460-LSmitll_SPLITT-OUT-X17-LSmitll_NOTT-INt X460-LSmitll_SPLITT-OUT-X88-LSmitll_NOTT-INt LSmitll_SPLITT

t1469 X461-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-INt 0 X461-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1470 X461-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-INt 0 X461-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X461 X465-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-IN X461-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-INt X461-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-INt LSmitll_SPLITT

t1471 X462-LSmitll_SPLITT-OUT-X299-LSmitll_DFFT-INt 0 X462-LSmitll_SPLITT-OUT-X299-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1472 X462-LSmitll_SPLITT-OUT-X305-LSmitll_DFFT-INt 0 X462-LSmitll_SPLITT-OUT-X305-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
X462 X464-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-IN X462-LSmitll_SPLITT-OUT-X299-LSmitll_DFFT-INt X462-LSmitll_SPLITT-OUT-X305-LSmitll_DFFT-INt LSmitll_SPLITT

t1473 X463-LSmitll_SPLITT-OUT-X288-LSmitll_DFFT-INt 0 X463-LSmitll_SPLITT-OUT-X288-LSmitll_DFFT-IN 0 z0=5 td=2.8ps
t1474 X463-LSmitll_SPLITT-OUT-X307-LSmitll_DFFT-INt 0 X463-LSmitll_SPLITT-OUT-X307-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X463 X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-IN X463-LSmitll_SPLITT-OUT-X288-LSmitll_DFFT-INt X463-LSmitll_SPLITT-OUT-X307-LSmitll_DFFT-INt LSmitll_SPLITT

t1475 X464-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-INt 0 X464-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1476 X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-INt 0 X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X464 X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-IN X464-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-INt X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-INt LSmitll_SPLITT

t1477 X465-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-INt 0 X465-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1478 X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-INt 0 X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X465 X472-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-IN X465-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-INt X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-INt LSmitll_SPLITT

t1479 X466-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-INt 0 X466-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
t1480 X466-LSmitll_SPLITT-OUT-X309-LSmitll_DFFT-INt 0 X466-LSmitll_SPLITT-OUT-X309-LSmitll_DFFT-IN 0 z0=5 td=3.0ps
X466 X468-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-IN X466-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-INt X466-LSmitll_SPLITT-OUT-X309-LSmitll_DFFT-INt LSmitll_SPLITT

t1481 X467-LSmitll_SPLITT-OUT-X11-LSmitll_DFFT-INt 0 X467-LSmitll_SPLITT-OUT-X11-LSmitll_DFFT-IN 0 z0=5 td=1.8ps
t1482 X467-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-INt 0 X467-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X467 X468-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-IN X467-LSmitll_SPLITT-OUT-X11-LSmitll_DFFT-INt X467-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-INt LSmitll_SPLITT

t1483 X468-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-INt 0 X468-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1484 X468-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-INt 0 X468-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X468 X471-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-IN X468-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-INt X468-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-INt LSmitll_SPLITT

t1485 X469-LSmitll_SPLITT-OUT-X306-LSmitll_DFFT-INt 0 X469-LSmitll_SPLITT-OUT-X306-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1486 X469-LSmitll_SPLITT-OUT-X311-LSmitll_OR2T-INt 0 X469-LSmitll_SPLITT-OUT-X311-LSmitll_OR2T-IN 0 z0=5 td=1.5ps
X469 X470-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-IN X469-LSmitll_SPLITT-OUT-X306-LSmitll_DFFT-INt X469-LSmitll_SPLITT-OUT-X311-LSmitll_OR2T-INt LSmitll_SPLITT

t1487 X470-LSmitll_SPLITT-OUT-X566-LSmitll_SPLITT-INt 0 X470-LSmitll_SPLITT-OUT-X566-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1488 X470-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-INt 0 X470-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X470 X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-IN X470-LSmitll_SPLITT-OUT-X566-LSmitll_SPLITT-INt X470-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-INt LSmitll_SPLITT

t1489 X471-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-INt 0 X471-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1490 X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-INt 0 X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
X471 X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-IN X471-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-INt X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-INt LSmitll_SPLITT

t1491 X472-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-INt 0 X472-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1492 X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-INt 0 X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X472 X486-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-IN X472-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-INt X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-INt LSmitll_SPLITT

t1493 X473-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-INt 0 X473-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-IN 0 z0=5 td=0.4ps
t1494 X473-LSmitll_SPLITT-OUT-X272-LSmitll_DFFT-INt 0 X473-LSmitll_SPLITT-OUT-X272-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
X473 X475-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-IN X473-LSmitll_SPLITT-OUT-X121-LSmitll_AND2T-INt X473-LSmitll_SPLITT-OUT-X272-LSmitll_DFFT-INt LSmitll_SPLITT

t1495 X474-LSmitll_SPLITT-OUT-X5-LSmitll_DFFT-INt 0 X474-LSmitll_SPLITT-OUT-X5-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
t1496 X474-LSmitll_SPLITT-OUT-X151-LSmitll_DFFT-INt 0 X474-LSmitll_SPLITT-OUT-X151-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
X474 X475-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-IN X474-LSmitll_SPLITT-OUT-X5-LSmitll_DFFT-INt X474-LSmitll_SPLITT-OUT-X151-LSmitll_DFFT-INt LSmitll_SPLITT

t1497 X475-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-INt 0 X475-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-IN 0 z0=5 td=0.6ps
t1498 X475-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-INt 0 X475-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X475 X478-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-IN X475-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-INt X475-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-INt LSmitll_SPLITT

t1499 X476-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-INt 0 X476-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
t1500 X476-LSmitll_SPLITT-OUT-X235-LSmitll_DFFT-INt 0 X476-LSmitll_SPLITT-OUT-X235-LSmitll_DFFT-IN 0 z0=5 td=3.6ps
X476 X477-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-IN X476-LSmitll_SPLITT-OUT-X26-LSmitll_AND2T-INt X476-LSmitll_SPLITT-OUT-X235-LSmitll_DFFT-INt LSmitll_SPLITT

t1501 X477-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-INt 0 X477-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1502 X477-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-INt 0 X477-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X477 X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-IN X477-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-INt X477-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-INt LSmitll_SPLITT

t1503 X478-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-INt 0 X478-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1504 X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-INt 0 X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X478 X485-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-IN X478-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-INt X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-INt LSmitll_SPLITT

t1505 X479-LSmitll_SPLITT-OUT-X169-LSmitll_DFFT-INt 0 X479-LSmitll_SPLITT-OUT-X169-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
t1506 X479-LSmitll_SPLITT-OUT-X300-LSmitll_DFFT-INt 0 X479-LSmitll_SPLITT-OUT-X300-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X479 X481-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-IN X479-LSmitll_SPLITT-OUT-X169-LSmitll_DFFT-INt X479-LSmitll_SPLITT-OUT-X300-LSmitll_DFFT-INt LSmitll_SPLITT

t1507 X480-LSmitll_SPLITT-OUT-X310-LSmitll_DFFT-INt 0 X480-LSmitll_SPLITT-OUT-X310-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1508 X480-LSmitll_SPLITT-OUT-X312-LSmitll_OR2T-INt 0 X480-LSmitll_SPLITT-OUT-X312-LSmitll_OR2T-IN 0 z0=5 td=0.5ps
X480 X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-IN X480-LSmitll_SPLITT-OUT-X310-LSmitll_DFFT-INt X480-LSmitll_SPLITT-OUT-X312-LSmitll_OR2T-INt LSmitll_SPLITT

t1509 X481-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-INt 0 X481-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1510 X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-INt 0 X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X481 X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-IN X481-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-INt X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-INt LSmitll_SPLITT

t1511 X482-LSmitll_SPLITT-OUT-X6-LSmitll_NOTT-INt 0 X482-LSmitll_SPLITT-OUT-X6-LSmitll_NOTT-IN 0 z0=5 td=0.7ps
t1512 X482-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-INt 0 X482-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-IN 0 z0=5 td=2.7ps
X482 X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-IN X482-LSmitll_SPLITT-OUT-X6-LSmitll_NOTT-INt X482-LSmitll_SPLITT-OUT-X24-LSmitll_AND2T-INt LSmitll_SPLITT

t1513 X483-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-INt 0 X483-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1514 X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-INt 0 X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X483 X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-IN X483-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-INt X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-INt LSmitll_SPLITT

t1515 X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-INt 0 X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1516 X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-INt 0 X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X484 X485-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-IN X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-INt X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-INt LSmitll_SPLITT

t1517 X485-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-INt 0 X485-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1518 X485-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-INt 0 X485-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X485 X486-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-IN X485-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-INt X485-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-INt LSmitll_SPLITT

t1519 X486-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-INt 0 X486-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-IN 0 z0=5 td=5.1ps
t1520 X486-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-INt 0 X486-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
X486 X487-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-IN X486-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-INt X486-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-INt LSmitll_SPLITT

t1521 X487-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-INt 0 X487-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
t1522 X487-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-INt 0 X487-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-IN 0 z0=5 td=3.6ps
X487 X545-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-IN X487-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-INt X487-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-INt LSmitll_SPLITT

t1523 X488-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-INt 0 X488-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-IN 0 z0=5 td=3.6ps
t1524 X488-LSmitll_SPLITT-OUT-X210-LSmitll_DFFT-INt 0 X488-LSmitll_SPLITT-OUT-X210-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
X488 X490-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-IN X488-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-INt X488-LSmitll_SPLITT-OUT-X210-LSmitll_DFFT-INt LSmitll_SPLITT

t1525 X489-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-INt 0 X489-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-IN 0 z0=5 td=2.0ps
t1526 X489-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-INt 0 X489-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
X489 X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-IN X489-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-INt X489-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-INt LSmitll_SPLITT

t1527 X490-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-INt 0 X490-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
t1528 X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-INt 0 X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X490 X494-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-IN X490-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-INt X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-INt LSmitll_SPLITT

t1529 X491-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-INt 0 X491-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-IN 0 z0=5 td=1.4ps
t1530 X491-LSmitll_SPLITT-OUT-X222-LSmitll_DFFT-INt 0 X491-LSmitll_SPLITT-OUT-X222-LSmitll_DFFT-IN 0 z0=5 td=3.7ps
X491 X493-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-IN X491-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-INt X491-LSmitll_SPLITT-OUT-X222-LSmitll_DFFT-INt LSmitll_SPLITT

t1531 X492-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-INt 0 X492-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t1532 X492-LSmitll_SPLITT-OUT-X204-LSmitll_DFFT-INt 0 X492-LSmitll_SPLITT-OUT-X204-LSmitll_DFFT-IN 0 z0=5 td=2.7ps
X492 X493-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-IN X492-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-INt X492-LSmitll_SPLITT-OUT-X204-LSmitll_DFFT-INt LSmitll_SPLITT

t1533 X493-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-INt 0 X493-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1534 X493-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-INt 0 X493-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X493 X494-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-IN X493-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-INt X493-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-INt LSmitll_SPLITT

t1535 X494-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-INt 0 X494-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-IN 0 z0=5 td=0.5ps
t1536 X494-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-INt 0 X494-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X494 X501-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-IN X494-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-INt X494-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-INt LSmitll_SPLITT

t1537 X495-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-INt 0 X495-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1538 X495-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-INt 0 X495-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-IN 0 z0=5 td=2.5ps
X495 X497-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-IN X495-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-INt X495-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-INt LSmitll_SPLITT

t1539 X496-LSmitll_SPLITT-OUT-X255-LSmitll_DFFT-INt 0 X496-LSmitll_SPLITT-OUT-X255-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1540 X496-LSmitll_SPLITT-OUT-X270-LSmitll_DFFT-INt 0 X496-LSmitll_SPLITT-OUT-X270-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
X496 X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-IN X496-LSmitll_SPLITT-OUT-X255-LSmitll_DFFT-INt X496-LSmitll_SPLITT-OUT-X270-LSmitll_DFFT-INt LSmitll_SPLITT

t1541 X497-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-INt 0 X497-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1542 X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-INt 0 X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X497 X500-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-IN X497-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-INt X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-INt LSmitll_SPLITT

t1543 X498-LSmitll_SPLITT-OUT-X193-LSmitll_DFFT-INt 0 X498-LSmitll_SPLITT-OUT-X193-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
t1544 X498-LSmitll_SPLITT-OUT-X221-LSmitll_DFFT-INt 0 X498-LSmitll_SPLITT-OUT-X221-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
X498 X499-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-IN X498-LSmitll_SPLITT-OUT-X193-LSmitll_DFFT-INt X498-LSmitll_SPLITT-OUT-X221-LSmitll_DFFT-INt LSmitll_SPLITT

t1545 X499-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-INt 0 X499-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1546 X499-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-INt 0 X499-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X499 X500-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-IN X499-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-INt X499-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-INt LSmitll_SPLITT

t1547 X500-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-INt 0 X500-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1548 X500-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-INt 0 X500-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-IN 0 z0=5 td=2.8ps
X500 X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-IN X500-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-INt X500-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-INt LSmitll_SPLITT

t1549 X501-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-INt 0 X501-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t1550 X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-INt 0 X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X501 X515-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-IN X501-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-INt X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-INt LSmitll_SPLITT

t1551 X502-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt 0 X502-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
t1552 X502-LSmitll_SPLITT-OUT-X238-LSmitll_OR2T-INt 0 X502-LSmitll_SPLITT-OUT-X238-LSmitll_OR2T-IN 0 z0=5 td=2.1ps
X502 X504-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-IN X502-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt X502-LSmitll_SPLITT-OUT-X238-LSmitll_OR2T-INt LSmitll_SPLITT

t1553 X503-LSmitll_SPLITT-OUT-X81-LSmitll_DFFT-INt 0 X503-LSmitll_SPLITT-OUT-X81-LSmitll_DFFT-IN 0 z0=5 td=3.2ps
t1554 X503-LSmitll_SPLITT-OUT-X280-LSmitll_NDROT-INt 0 X503-LSmitll_SPLITT-OUT-X280-LSmitll_NDROT-IN 0 z0=5 td=3.0ps
X503 X504-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-IN X503-LSmitll_SPLITT-OUT-X81-LSmitll_DFFT-INt X503-LSmitll_SPLITT-OUT-X280-LSmitll_NDROT-INt LSmitll_SPLITT

t1555 X504-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-INt 0 X504-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1556 X504-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-INt 0 X504-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X504 X507-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-IN X504-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-INt X504-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-INt LSmitll_SPLITT

t1557 X505-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-INt 0 X505-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t1558 X505-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-INt 0 X505-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
X505 X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-IN X505-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-INt X505-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-INt LSmitll_SPLITT

t1559 X506-LSmitll_SPLITT-OUT-X564-LSmitll_SPLITT-INt 0 X506-LSmitll_SPLITT-OUT-X564-LSmitll_SPLITT-IN 0 z0=5 td=3.2ps
t1560 X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-INt 0 X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X506 X507-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-IN X506-LSmitll_SPLITT-OUT-X564-LSmitll_SPLITT-INt X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-INt LSmitll_SPLITT

t1561 X507-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-INt 0 X507-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1562 X507-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-INt 0 X507-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X507 X514-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-IN X507-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-INt X507-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-INt LSmitll_SPLITT

t1563 X508-LSmitll_SPLITT-OUT-X131-LSmitll_AND2T-INt 0 X508-LSmitll_SPLITT-OUT-X131-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
t1564 X508-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt 0 X508-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN 0 z0=5 td=2.8ps
X508 X510-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-IN X508-LSmitll_SPLITT-OUT-X131-LSmitll_AND2T-INt X508-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt LSmitll_SPLITT

t1565 X509-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-INt 0 X509-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
t1566 X509-LSmitll_SPLITT-OUT-X154-LSmitll_OR2T-INt 0 X509-LSmitll_SPLITT-OUT-X154-LSmitll_OR2T-IN 0 z0=5 td=1.0ps
X509 X510-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-IN X509-LSmitll_SPLITT-OUT-X133-LSmitll_AND2T-INt X509-LSmitll_SPLITT-OUT-X154-LSmitll_OR2T-INt LSmitll_SPLITT

t1567 X510-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-INt 0 X510-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1568 X510-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-INt 0 X510-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X510 X513-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-IN X510-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-INt X510-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-INt LSmitll_SPLITT

t1569 X511-LSmitll_SPLITT-OUT-X189-LSmitll_DFFT-INt 0 X511-LSmitll_SPLITT-OUT-X189-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
t1570 X511-LSmitll_SPLITT-OUT-X291-LSmitll_DFFT-INt 0 X511-LSmitll_SPLITT-OUT-X291-LSmitll_DFFT-IN 0 z0=5 td=3.6ps
X511 X512-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-IN X511-LSmitll_SPLITT-OUT-X189-LSmitll_DFFT-INt X511-LSmitll_SPLITT-OUT-X291-LSmitll_DFFT-INt LSmitll_SPLITT

t1571 X512-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-INt 0 X512-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1572 X512-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-INt 0 X512-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X512 X513-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-IN X512-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-INt X512-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-INt LSmitll_SPLITT

t1573 X513-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-INt 0 X513-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1574 X513-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-INt 0 X513-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X513 X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-IN X513-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-INt X513-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-INt LSmitll_SPLITT

t1575 X514-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-INt 0 X514-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1576 X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-INt 0 X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X514 X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-IN X514-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-INt X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-INt LSmitll_SPLITT

t1577 X515-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-INt 0 X515-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-IN 0 z0=5 td=3.5ps
t1578 X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-INt 0 X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-IN 0 z0=5 td=5.0ps
X515 X544-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-IN X515-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-INt X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-INt LSmitll_SPLITT

t1579 X516-LSmitll_SPLITT-OUT-X198-LSmitll_DFFT-INt 0 X516-LSmitll_SPLITT-OUT-X198-LSmitll_DFFT-IN 0 z0=5 td=0.4ps
t1580 X516-LSmitll_SPLITT-OUT-X247-LSmitll_DFFT-INt 0 X516-LSmitll_SPLITT-OUT-X247-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X516 X518-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-IN X516-LSmitll_SPLITT-OUT-X198-LSmitll_DFFT-INt X516-LSmitll_SPLITT-OUT-X247-LSmitll_DFFT-INt LSmitll_SPLITT

t1581 X517-LSmitll_SPLITT-OUT-X223-LSmitll_DFFT-INt 0 X517-LSmitll_SPLITT-OUT-X223-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
t1582 X517-LSmitll_SPLITT-OUT-X286-LSmitll_DFFT-INt 0 X517-LSmitll_SPLITT-OUT-X286-LSmitll_DFFT-IN 0 z0=5 td=2.0ps
X517 X518-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-IN X517-LSmitll_SPLITT-OUT-X223-LSmitll_DFFT-INt X517-LSmitll_SPLITT-OUT-X286-LSmitll_DFFT-INt LSmitll_SPLITT

t1583 X518-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-INt 0 X518-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1584 X518-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-INt 0 X518-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-IN 0 z0=5 td=1.0ps
X518 X522-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-IN X518-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-INt X518-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-INt LSmitll_SPLITT

t1585 X519-LSmitll_SPLITT-OUT-X155-LSmitll_OR2T-INt 0 X519-LSmitll_SPLITT-OUT-X155-LSmitll_OR2T-IN 0 z0=5 td=1.4ps
t1586 X519-LSmitll_SPLITT-OUT-X162-LSmitll_DFFT-INt 0 X519-LSmitll_SPLITT-OUT-X162-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X519 X521-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-IN X519-LSmitll_SPLITT-OUT-X155-LSmitll_OR2T-INt X519-LSmitll_SPLITT-OUT-X162-LSmitll_DFFT-INt LSmitll_SPLITT

t1587 X520-LSmitll_SPLITT-OUT-X206-LSmitll_DFFT-INt 0 X520-LSmitll_SPLITT-OUT-X206-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
t1588 X520-LSmitll_SPLITT-OUT-X234-LSmitll_DFFT-INt 0 X520-LSmitll_SPLITT-OUT-X234-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
X520 X521-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-IN X520-LSmitll_SPLITT-OUT-X206-LSmitll_DFFT-INt X520-LSmitll_SPLITT-OUT-X234-LSmitll_DFFT-INt LSmitll_SPLITT

t1589 X521-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-INt 0 X521-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t1590 X521-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-INt 0 X521-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X521 X522-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-IN X521-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-INt X521-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-INt LSmitll_SPLITT

t1591 X522-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-INt 0 X522-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-IN 0 z0=5 td=4.2ps
t1592 X522-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-INt 0 X522-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
X522 X529-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-IN X522-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-INt X522-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-INt LSmitll_SPLITT

t1593 X523-LSmitll_SPLITT-OUT-X211-LSmitll_DFFT-INt 0 X523-LSmitll_SPLITT-OUT-X211-LSmitll_DFFT-IN 0 z0=5 td=1.7ps
t1594 X523-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-INt 0 X523-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
X523 X525-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-IN X523-LSmitll_SPLITT-OUT-X211-LSmitll_DFFT-INt X523-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-INt LSmitll_SPLITT

t1595 X524-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-INt 0 X524-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t1596 X524-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-INt 0 X524-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
X524 X525-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-IN X524-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-INt X524-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-INt LSmitll_SPLITT

t1597 X525-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-INt 0 X525-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
t1598 X525-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-INt 0 X525-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
X525 X528-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-IN X525-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-INt X525-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-INt LSmitll_SPLITT

t1599 X526-LSmitll_SPLITT-OUT-X246-LSmitll_DFFT-INt 0 X526-LSmitll_SPLITT-OUT-X246-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
t1600 X526-LSmitll_SPLITT-OUT-X254-LSmitll_DFFT-INt 0 X526-LSmitll_SPLITT-OUT-X254-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X526 X527-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-IN X526-LSmitll_SPLITT-OUT-X246-LSmitll_DFFT-INt X526-LSmitll_SPLITT-OUT-X254-LSmitll_DFFT-INt LSmitll_SPLITT

t1601 X527-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-INt 0 X527-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1602 X527-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-INt 0 X527-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X527 X528-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-IN X527-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-INt X527-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-INt LSmitll_SPLITT

t1603 X528-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-INt 0 X528-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t1604 X528-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-INt 0 X528-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X528 X529-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-IN X528-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-INt X528-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-INt LSmitll_SPLITT

t1605 X529-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-INt 0 X529-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1606 X529-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-INt 0 X529-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X529 X543-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-IN X529-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-INt X529-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-INt LSmitll_SPLITT

t1607 X530-LSmitll_SPLITT-OUT-X85-LSmitll_DFFT-INt 0 X530-LSmitll_SPLITT-OUT-X85-LSmitll_DFFT-IN 0 z0=5 td=3.5ps
t1608 X530-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-INt 0 X530-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X530 X532-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-IN X530-LSmitll_SPLITT-OUT-X85-LSmitll_DFFT-INt X530-LSmitll_SPLITT-OUT-X251-LSmitll_AND2T-INt LSmitll_SPLITT

t1609 X531-LSmitll_SPLITT-OUT-X86-LSmitll_DFFT-INt 0 X531-LSmitll_SPLITT-OUT-X86-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1610 X531-LSmitll_SPLITT-OUT-X134-LSmitll_AND2T-INt 0 X531-LSmitll_SPLITT-OUT-X134-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X531 X532-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-IN X531-LSmitll_SPLITT-OUT-X86-LSmitll_DFFT-INt X531-LSmitll_SPLITT-OUT-X134-LSmitll_AND2T-INt LSmitll_SPLITT

t1611 X532-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-INt 0 X532-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
t1612 X532-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-INt 0 X532-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X532 X535-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-IN X532-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-INt X532-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-INt LSmitll_SPLITT

t1613 X533-LSmitll_SPLITT-OUT-X173-LSmitll_DFFT-INt 0 X533-LSmitll_SPLITT-OUT-X173-LSmitll_DFFT-IN 0 z0=5 td=1.7ps
t1614 X533-LSmitll_SPLITT-OUT-X174-LSmitll_DFFT-INt 0 X533-LSmitll_SPLITT-OUT-X174-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
X533 X534-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-IN X533-LSmitll_SPLITT-OUT-X173-LSmitll_DFFT-INt X533-LSmitll_SPLITT-OUT-X174-LSmitll_DFFT-INt LSmitll_SPLITT

t1615 X534-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-INt 0 X534-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-IN 0 z0=5 td=11.7ps
t1616 X534-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-INt 0 X534-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X534 X535-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-IN X534-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-INt X534-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-INt LSmitll_SPLITT

t1617 X535-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-INt 0 X535-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1618 X535-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-INt 0 X535-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X535 X542-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-IN X535-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-INt X535-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-INt LSmitll_SPLITT

t1619 X536-LSmitll_SPLITT-OUT-X269-LSmitll_DFFT-INt 0 X536-LSmitll_SPLITT-OUT-X269-LSmitll_DFFT-IN 0 z0=5 td=3.8ps
t1620 X536-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-INt 0 X536-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X536 X538-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-IN X536-LSmitll_SPLITT-OUT-X269-LSmitll_DFFT-INt X536-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-INt LSmitll_SPLITT

t1621 X537-LSmitll_SPLITT-OUT-X260-LSmitll_DFFT-INt 0 X537-LSmitll_SPLITT-OUT-X260-LSmitll_DFFT-IN 0 z0=5 td=3.1ps
t1622 X537-LSmitll_SPLITT-OUT-X302-LSmitll_DFFT-INt 0 X537-LSmitll_SPLITT-OUT-X302-LSmitll_DFFT-IN 0 z0=5 td=2.5ps
X537 X538-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-IN X537-LSmitll_SPLITT-OUT-X260-LSmitll_DFFT-INt X537-LSmitll_SPLITT-OUT-X302-LSmitll_DFFT-INt LSmitll_SPLITT

t1623 X538-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-INt 0 X538-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1624 X538-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-INt 0 X538-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X538 X541-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-IN X538-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-INt X538-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-INt LSmitll_SPLITT

t1625 X539-LSmitll_SPLITT-OUT-X172-LSmitll_DFFT-INt 0 X539-LSmitll_SPLITT-OUT-X172-LSmitll_DFFT-IN 0 z0=5 td=2.0ps
t1626 X539-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-INt 0 X539-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X539 X540-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-IN X539-LSmitll_SPLITT-OUT-X172-LSmitll_DFFT-INt X539-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-INt LSmitll_SPLITT

t1627 X540-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-INt 0 X540-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1628 X540-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-INt 0 X540-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X540 X541-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-IN X540-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-INt X540-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-INt LSmitll_SPLITT

t1629 X541-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-INt 0 X541-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
t1630 X541-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-INt 0 X541-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X541 X542-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-IN X541-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-INt X541-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-INt LSmitll_SPLITT

t1631 X542-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-INt 0 X542-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
t1632 X542-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-INt 0 X542-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
X542 X543-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-IN X542-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-INt X542-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-INt LSmitll_SPLITT

t1633 X543-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-INt 0 X543-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-IN 0 z0=5 td=5.9ps
t1634 X543-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-INt 0 X543-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-IN 0 z0=5 td=6.6ps
X543 X544-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-IN X543-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-INt X543-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-INt LSmitll_SPLITT

t1635 X544-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-INt 0 X544-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-IN 0 z0=5 td=4.0ps
t1636 X544-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-INt 0 X544-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-IN 0 z0=5 td=5.3ps
X544 X545-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-IN X544-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-INt X544-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-INt LSmitll_SPLITT

t1637 X545-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-INt 0 X545-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-IN 0 z0=5 td=7.6ps
t1638 X545-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-INt 0 X545-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-IN 0 z0=5 td=5.5ps
X545 X567-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-IN X545-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-INt X545-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-INt LSmitll_SPLITT

t1639 X546-LSmitll_SPLITT-OUT-X4-LSmitll_NOTT-INt 0 X546-LSmitll_SPLITT-OUT-X4-LSmitll_NOTT-IN 0 z0=5 td=0.7ps
t1640 X546-SPLITT-OUT-R-INt 0 X546-SPLITT-OUT-R-IN 0 z0=5 td=10.1ps
X546 X483-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-IN X546-LSmitll_SPLITT-OUT-X4-LSmitll_NOTT-INt X546-SPLITT-OUT-R-INt LSmitll_SPLITT

t1641 X547-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-INt 0 X547-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-IN 0 z0=5 td=0.7ps
t1642 X547-SPLITT-OUT-R-INt 0 X547-SPLITT-OUT-R-IN 0 z0=5 td=5.0ps
X547 X477-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-IN X547-LSmitll_SPLITT-OUT-X25-LSmitll_AND2T-INt X547-SPLITT-OUT-R-INt LSmitll_SPLITT

t1643 X548-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-INt 0 X548-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1644 X548-SPLITT-OUT-R-INt 0 X548-SPLITT-OUT-R-IN 0 z0=5 td=4.8ps
X548 X353-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-IN X548-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-INt X548-SPLITT-OUT-R-INt LSmitll_SPLITT

t1645 X549-LSmitll_SPLITT-OUT-X68-LSmitll_DFFT-INt 0 X549-LSmitll_SPLITT-OUT-X68-LSmitll_DFFT-IN 0 z0=5 td=0.4ps
t1646 X549-SPLITT-OUT-R-INt 0 X549-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X549 X360-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-IN X549-LSmitll_SPLITT-OUT-X68-LSmitll_DFFT-INt X549-SPLITT-OUT-R-INt LSmitll_SPLITT

t1647 X550-LSmitll_SPLITT-OUT-X82-LSmitll_DFFT-INt 0 X550-LSmitll_SPLITT-OUT-X82-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1648 X550-SPLITT-OUT-R-INt 0 X550-SPLITT-OUT-R-IN 0 z0=5 td=4.3ps
X550 X411-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-IN X550-LSmitll_SPLITT-OUT-X82-LSmitll_DFFT-INt X550-SPLITT-OUT-R-INt LSmitll_SPLITT

t1649 X551-LSmitll_SPLITT-OUT-X116-LSmitll_DFFT-INt 0 X551-LSmitll_SPLITT-OUT-X116-LSmitll_DFFT-IN 0 z0=5 td=0.4ps
t1650 X551-SPLITT-OUT-R-INt 0 X551-SPLITT-OUT-R-IN 0 z0=5 td=5.2ps
X551 X366-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-IN X551-LSmitll_SPLITT-OUT-X116-LSmitll_DFFT-INt X551-SPLITT-OUT-R-INt LSmitll_SPLITT

t1651 X552-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt 0 X552-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN 0 z0=5 td=0.7ps
t1652 X552-SPLITT-OUT-R-INt 0 X552-SPLITT-OUT-R-IN 0 z0=5 td=7.1ps
X552 X338-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-IN X552-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt X552-SPLITT-OUT-R-INt LSmitll_SPLITT

t1653 X553-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-INt 0 X553-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1654 X553-SPLITT-OUT-R-INt 0 X553-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X553 X499-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-IN X553-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-INt X553-SPLITT-OUT-R-INt LSmitll_SPLITT

t1655 X554-LSmitll_SPLITT-OUT-X175-LSmitll_DFFT-INt 0 X554-LSmitll_SPLITT-OUT-X175-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1656 X554-SPLITT-OUT-R-INt 0 X554-SPLITT-OUT-R-IN 0 z0=5 td=9.7ps
X554 X382-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-IN X554-LSmitll_SPLITT-OUT-X175-LSmitll_DFFT-INt X554-SPLITT-OUT-R-INt LSmitll_SPLITT

t1657 X555-LSmitll_SPLITT-OUT-X182-LSmitll_DFFT-INt 0 X555-LSmitll_SPLITT-OUT-X182-LSmitll_DFFT-IN 0 z0=5 td=0.4ps
t1658 X555-SPLITT-OUT-R-INt 0 X555-SPLITT-OUT-R-IN 0 z0=5 td=3.3ps
X555 X455-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-IN X555-LSmitll_SPLITT-OUT-X182-LSmitll_DFFT-INt X555-SPLITT-OUT-R-INt LSmitll_SPLITT

t1659 X556-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-INt 0 X556-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1660 X556-SPLITT-OUT-R-INt 0 X556-SPLITT-OUT-R-IN 0 z0=5 td=10.0ps
X556 X540-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-IN X556-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-INt X556-SPLITT-OUT-R-INt LSmitll_SPLITT

t1661 X557-LSmitll_SPLITT-OUT-X190-LSmitll_DFFT-INt 0 X557-LSmitll_SPLITT-OUT-X190-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1662 X557-SPLITT-OUT-R-INt 0 X557-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X557 X512-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-IN X557-LSmitll_SPLITT-OUT-X190-LSmitll_DFFT-INt X557-SPLITT-OUT-R-INt LSmitll_SPLITT

t1663 X558-LSmitll_SPLITT-OUT-X236-LSmitll_DFFT-INt 0 X558-LSmitll_SPLITT-OUT-X236-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1664 X558-SPLITT-OUT-R-INt 0 X558-SPLITT-OUT-R-IN 0 z0=5 td=4.8ps
X558 X324-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-IN X558-LSmitll_SPLITT-OUT-X236-LSmitll_DFFT-INt X558-SPLITT-OUT-R-INt LSmitll_SPLITT

t1665 X559-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-INt 0 X559-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-IN 0 z0=5 td=0.8ps
t1666 X559-SPLITT-OUT-R-INt 0 X559-SPLITT-OUT-R-IN 0 z0=5 td=3.7ps
X559 X534-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-IN X559-LSmitll_SPLITT-OUT-X250-LSmitll_XORT-INt X559-SPLITT-OUT-R-INt LSmitll_SPLITT

t1667 X560-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-INt 0 X560-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1668 X560-SPLITT-OUT-R-INt 0 X560-SPLITT-OUT-R-IN 0 z0=5 td=4.3ps
X560 X396-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-IN X560-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-INt X560-SPLITT-OUT-R-INt LSmitll_SPLITT

t1669 X561-LSmitll_SPLITT-OUT-X285-LSmitll_DFFT-INt 0 X561-LSmitll_SPLITT-OUT-X285-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1670 X561-SPLITT-OUT-R-INt 0 X561-SPLITT-OUT-R-IN 0 z0=5 td=9.9ps
X561 X527-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-IN X561-LSmitll_SPLITT-OUT-X285-LSmitll_DFFT-INt X561-SPLITT-OUT-R-INt LSmitll_SPLITT

t1671 X562-LSmitll_SPLITT-OUT-X287-LSmitll_DFFT-INt 0 X562-LSmitll_SPLITT-OUT-X287-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1672 X562-SPLITT-OUT-R-INt 0 X562-SPLITT-OUT-R-IN 0 z0=5 td=3.3ps
X562 X441-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-IN X562-LSmitll_SPLITT-OUT-X287-LSmitll_DFFT-INt X562-SPLITT-OUT-R-INt LSmitll_SPLITT

t1673 X563-LSmitll_SPLITT-OUT-X292-LSmitll_DFFT-INt 0 X563-LSmitll_SPLITT-OUT-X292-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1674 X563-SPLITT-OUT-R-INt 0 X563-SPLITT-OUT-R-IN 0 z0=5 td=4.7ps
X563 X418-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-IN X563-LSmitll_SPLITT-OUT-X292-LSmitll_DFFT-INt X563-SPLITT-OUT-R-INt LSmitll_SPLITT

t1675 X564-LSmitll_SPLITT-OUT-X293-LSmitll_NOTT-INt 0 X564-LSmitll_SPLITT-OUT-X293-LSmitll_NOTT-IN 0 z0=5 td=0.7ps
t1676 X564-SPLITT-OUT-R-INt 0 X564-SPLITT-OUT-R-IN 0 z0=5 td=9.7ps
X564 X506-LSmitll_SPLITT-OUT-X564-LSmitll_SPLITT-IN X564-LSmitll_SPLITT-OUT-X293-LSmitll_NOTT-INt X564-SPLITT-OUT-R-INt LSmitll_SPLITT

t1677 X565-LSmitll_SPLITT-OUT-X294-LSmitll_NOTT-INt 0 X565-LSmitll_SPLITT-OUT-X294-LSmitll_NOTT-IN 0 z0=5 td=0.7ps
t1678 X565-SPLITT-OUT-R-INt 0 X565-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X565 X424-LSmitll_SPLITT-OUT-X565-LSmitll_SPLITT-IN X565-LSmitll_SPLITT-OUT-X294-LSmitll_NOTT-INt X565-SPLITT-OUT-R-INt LSmitll_SPLITT

t1679 X566-LSmitll_SPLITT-OUT-X308-LSmitll_DFFT-INt 0 X566-LSmitll_SPLITT-OUT-X308-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1680 X566-SPLITT-OUT-R-INt 0 X566-SPLITT-OUT-R-IN 0 z0=5 td=7.4ps
X566 X470-LSmitll_SPLITT-OUT-X566-LSmitll_SPLITT-IN X566-LSmitll_SPLITT-OUT-X308-LSmitll_DFFT-INt X566-SPLITT-OUT-R-INt LSmitll_SPLITT

t1681 X567-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-INt 0 X567-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-IN 0 z0=5 td=8.3ps
t1682 X567-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-INt 0 X567-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-IN 0 z0=5 td=6.4ps
X567 GCLK X567-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-INt X567-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-INt LSmitll_SPLITT

* PTLs from input pads
t783 GCLKt 0 GCLK 0 z0=5 td=13.1ps
t571 bit7t 0 bit7 0 z0=5 td=16.3ps
t575 bit6t 0 bit6 0 z0=5 td=15.7ps
t579 bit5t 0 bit5 0 z0=5 td=9.9ps
t583 bit4t 0 bit4 0 z0=5 td=11.9ps
t587 bit3t 0 bit3 0 z0=5 td=12.3ps
t591 bit2t 0 bit2 0 z0=5 td=10.1ps
t595 bit1t 0 bit1 0 z0=5 td=9.2ps

t599 overflowt 0 overflow 0 z0=5 td=9.3ps
t603 zerot 0 zero 0 z0=5 td=6.3ps
t607 negt 0 neg 0 z0=5 td=7.9ps

* PTLs to output pads
t961 Imm0t 0 Imm0 0 z0=5 td=8.4ps
t964 Imm1t 0 Imm1 0 z0=5 td=13.9ps
t967 Imm2t 0 Imm2 0 z0=5 td=15.0ps
t970 Imm3t 0 Imm3 0 z0=5 td=6.5ps
t1164 select0t 0 select0 0 z0=5 td=3.9ps
t1163 select1t 0 select1 0 z0=5 td=2.8ps
t953 readt 0 read 0 z0=5 td=13.3ps
t1171 Addr0t 0 Addr0 0 z0=5 td=3.3ps
t1172 Addr1t 0 Addr1 0 z0=5 td=3.5ps
t1162 write_flagst 0 write_flags 0 z0=5 td=3.1ps

t1023 Op_Aritht 0 Op_Arith 0 z0=5 td=5.5ps
t1024 Op_Andt 0 Op_And 0 z0=5 td=5.9ps
t1025 Op_Xort 0 Op_Xor 0 z0=5 td=2.6ps
t1026 Cmpl_b0t 0 Cmpl_b0 0 z0=5 td=5.9ps
t1027 Cmpl_b1t 0 Cmpl_b1 0 z0=5 td=4.4ps
t1028 Cint 0 Cin 0 z0=5 td=3.5ps

t1130 readNextInstr0t 0 readNextInstr0 0 z0=5 td=4.9ps
t1131 readNextInstr1t 0 readNextInstr1 0 z0=5 td=8.9ps
t1126 nextInstrAddr0_0t 0 nextInstrAddr0_0 0 z0=5 td=4.2ps
t1127 nextInstrAddr0_1t 0 nextInstrAddr0_1 0 z0=5 td=3.8ps
t1128 nextInstrAddr1_0t 0 nextInstrAddr1_0 0 z0=5 td=5.4ps
t1129 nextInstrAddr1_1t 0 nextInstrAddr1_1 0 z0=5 td=5.3ps

.ends Control_Unit_final_route