.subckt ALU_Reg_file_final_route Imm3t Imm2t Imm1t Imm0t select1t select0t readt addr0t addr1t write_flagst Op_Aritht Op_Andt Op_Xort Cmpl_b1t Cmpl_b0t Cint GCLKt reg1_out0_pad reg1_out1_pad reg1_out2_pad reg1_out3_pad reg2_out0_pad reg2_out1_pad reg2_out2_pad reg2_out3_pad regFlags_out0 regFlags_out0_pad regFlags_out1 regFlags_out1_pad regFlags_out2 regFlags_out2_pad

X685 X519-SPLITT-OUT-R-IN X519-SPLITT-OUT-R-INr LSmitll_PTLRX
X686 X519-SPLITT-OUT-R-INr X519-SPLITT-OUT-R-INdc LSmitll_SFQDC
R687 X519-SPLITT-OUT-R-INdc 0 5
X688 X519-SPLITT-OUT-R-IN PAD

X689 X520-SPLITT-OUT-R-IN X520-SPLITT-OUT-R-INr LSmitll_PTLRX
X690 X520-SPLITT-OUT-R-INr X520-SPLITT-OUT-R-INdc LSmitll_SFQDC
R691 X520-SPLITT-OUT-R-INdc 0 5
X692 X520-SPLITT-OUT-R-IN PAD

X693 X521-SPLITT-OUT-R-IN X521-SPLITT-OUT-R-INr LSmitll_PTLRX
X694 X521-SPLITT-OUT-R-INr X521-SPLITT-OUT-R-INdc LSmitll_SFQDC
R695 X521-SPLITT-OUT-R-INdc 0 5
X696 X521-SPLITT-OUT-R-IN PAD

X697 X522-SPLITT-OUT-R-IN X522-SPLITT-OUT-R-INr LSmitll_PTLRX
X698 X522-SPLITT-OUT-R-INr X522-SPLITT-OUT-R-INdc LSmitll_SFQDC
R699 X522-SPLITT-OUT-R-INdc 0 5
X700 X522-SPLITT-OUT-R-IN PAD

X701 X523-SPLITT-OUT-R-IN X523-SPLITT-OUT-R-INr LSmitll_PTLRX
X702 X523-SPLITT-OUT-R-INr X523-SPLITT-OUT-R-INdc LSmitll_SFQDC
R703 X523-SPLITT-OUT-R-INdc 0 5
X704 X523-SPLITT-OUT-R-IN PAD

X705 X524-SPLITT-OUT-R-IN X524-SPLITT-OUT-R-INr LSmitll_PTLRX
X706 X524-SPLITT-OUT-R-INr X524-SPLITT-OUT-R-INdc LSmitll_SFQDC
R707 X524-SPLITT-OUT-R-INdc 0 5
X708 X524-SPLITT-OUT-R-IN PAD

X709 X525-SPLITT-OUT-R-IN X525-SPLITT-OUT-R-INr LSmitll_PTLRX
X710 X525-SPLITT-OUT-R-INr X525-SPLITT-OUT-R-INdc LSmitll_SFQDC
R711 X525-SPLITT-OUT-R-INdc 0 5
X712 X525-SPLITT-OUT-R-IN PAD

X713 X526-SPLITT-OUT-R-IN X526-SPLITT-OUT-R-INr LSmitll_PTLRX
X714 X526-SPLITT-OUT-R-INr X526-SPLITT-OUT-R-INdc LSmitll_SFQDC
R715 X526-SPLITT-OUT-R-INdc 0 5
X716 X526-SPLITT-OUT-R-IN PAD

X717 X527-SPLITT-OUT-R-IN X527-SPLITT-OUT-R-INr LSmitll_PTLRX
X718 X527-SPLITT-OUT-R-INr X527-SPLITT-OUT-R-INdc LSmitll_SFQDC
R719 X527-SPLITT-OUT-R-INdc 0 5
X720 X527-SPLITT-OUT-R-IN PAD

X721 X528-SPLITT-OUT-R-IN X528-SPLITT-OUT-R-INr LSmitll_PTLRX
X722 X528-SPLITT-OUT-R-INr X528-SPLITT-OUT-R-INdc LSmitll_SFQDC
R723 X528-SPLITT-OUT-R-INdc 0 5
X724 X528-SPLITT-OUT-R-IN PAD

X725 X529-SPLITT-OUT-R-IN X529-SPLITT-OUT-R-INr LSmitll_PTLRX
X726 X529-SPLITT-OUT-R-INr X529-SPLITT-OUT-R-INdc LSmitll_SFQDC
R727 X529-SPLITT-OUT-R-INdc 0 5
X728 X529-SPLITT-OUT-R-IN PAD

X729 X530-SPLITT-OUT-R-IN X530-SPLITT-OUT-R-INr LSmitll_PTLRX
X730 X530-SPLITT-OUT-R-INr X530-SPLITT-OUT-R-INdc LSmitll_SFQDC
R731 X530-SPLITT-OUT-R-INdc 0 5
X732 X530-SPLITT-OUT-R-IN PAD

X733 X531-SPLITT-OUT-R-IN X531-SPLITT-OUT-R-INr LSmitll_PTLRX
X734 X531-SPLITT-OUT-R-INr X531-SPLITT-OUT-R-INdc LSmitll_SFQDC
R735 X531-SPLITT-OUT-R-INdc 0 5
X736 X531-SPLITT-OUT-R-IN PAD

X737 X532-SPLITT-OUT-R-IN X532-SPLITT-OUT-R-INr LSmitll_PTLRX
X738 X532-SPLITT-OUT-R-INr X532-SPLITT-OUT-R-INdc LSmitll_SFQDC
R739 X532-SPLITT-OUT-R-INdc 0 5
X740 X532-SPLITT-OUT-R-IN PAD

X741 X533-SPLITT-OUT-R-IN X533-SPLITT-OUT-R-INr LSmitll_PTLRX
X742 X533-SPLITT-OUT-R-INr X533-SPLITT-OUT-R-INdc LSmitll_SFQDC
R743 X533-SPLITT-OUT-R-INdc 0 5
X744 X533-SPLITT-OUT-R-IN PAD

X745 X534-SPLITT-OUT-R-IN X534-SPLITT-OUT-R-INr LSmitll_PTLRX
X746 X534-SPLITT-OUT-R-INr X534-SPLITT-OUT-R-INdc LSmitll_SFQDC
R747 X534-SPLITT-OUT-R-INdc 0 5
X748 X534-SPLITT-OUT-R-IN PAD

X749 X535-SPLITT-OUT-R-IN X535-SPLITT-OUT-R-INr LSmitll_PTLRX
X750 X535-SPLITT-OUT-R-INr X535-SPLITT-OUT-R-INdc LSmitll_SFQDC
R751 X535-SPLITT-OUT-R-INdc 0 5
X752 X535-SPLITT-OUT-R-IN PAD

X753 X536-SPLITT-OUT-R-IN X536-SPLITT-OUT-R-INr LSmitll_PTLRX
X754 X536-SPLITT-OUT-R-INr X536-SPLITT-OUT-R-INdc LSmitll_SFQDC
R755 X536-SPLITT-OUT-R-INdc 0 5
X756 X536-SPLITT-OUT-R-IN PAD

X757 X537-SPLITT-OUT-R-IN X537-SPLITT-OUT-R-INr LSmitll_PTLRX
X758 X537-SPLITT-OUT-R-INr X537-SPLITT-OUT-R-INdc LSmitll_SFQDC
R759 X537-SPLITT-OUT-R-INdc 0 5
X760 X537-SPLITT-OUT-R-IN PAD

X761 X538-SPLITT-OUT-R-IN X538-SPLITT-OUT-R-INr LSmitll_PTLRX
X762 X538-SPLITT-OUT-R-INr X538-SPLITT-OUT-R-INdc LSmitll_SFQDC
R763 X538-SPLITT-OUT-R-INdc 0 5
X764 X538-SPLITT-OUT-R-IN PAD

X765 X539-SPLITT-OUT-R-IN X539-SPLITT-OUT-R-INr LSmitll_PTLRX
X766 X539-SPLITT-OUT-R-INr X539-SPLITT-OUT-R-INdc LSmitll_SFQDC
R767 X539-SPLITT-OUT-R-INdc 0 5
X768 X539-SPLITT-OUT-R-IN PAD

X769 X540-SPLITT-OUT-R-IN X540-SPLITT-OUT-R-INr LSmitll_PTLRX
X770 X540-SPLITT-OUT-R-INr X540-SPLITT-OUT-R-INdc LSmitll_SFQDC
R771 X540-SPLITT-OUT-R-INdc 0 5
X772 X540-SPLITT-OUT-R-IN PAD

X773 X541-SPLITT-OUT-R-IN X541-SPLITT-OUT-R-INr LSmitll_PTLRX
X774 X541-SPLITT-OUT-R-INr X541-SPLITT-OUT-R-INdc LSmitll_SFQDC
R775 X541-SPLITT-OUT-R-INdc 0 5
X776 X541-SPLITT-OUT-R-IN PAD

X777 X542-SPLITT-OUT-R-IN X542-SPLITT-OUT-R-INr LSmitll_PTLRX
X778 X542-SPLITT-OUT-R-INr X542-SPLITT-OUT-R-INdc LSmitll_SFQDC
R779 X542-SPLITT-OUT-R-INdc 0 5
X780 X542-SPLITT-OUT-R-IN PAD

X781 X543-SPLITT-OUT-R-IN X543-SPLITT-OUT-R-INr LSmitll_PTLRX
X782 X543-SPLITT-OUT-R-INr X543-SPLITT-OUT-R-INdc LSmitll_SFQDC
R783 X543-SPLITT-OUT-R-INdc 0 5
X784 X543-SPLITT-OUT-R-IN PAD

X785 X544-SPLITT-OUT-R-IN X544-SPLITT-OUT-R-INr LSmitll_PTLRX
X786 X544-SPLITT-OUT-R-INr X544-SPLITT-OUT-R-INdc LSmitll_SFQDC
R787 X544-SPLITT-OUT-R-INdc 0 5
X788 X544-SPLITT-OUT-R-IN PAD

X789 X545-SPLITT-OUT-R-IN X545-SPLITT-OUT-R-INr LSmitll_PTLRX
X790 X545-SPLITT-OUT-R-INr X545-SPLITT-OUT-R-INdc LSmitll_SFQDC
R791 X545-SPLITT-OUT-R-INdc 0 5
X792 X545-SPLITT-OUT-R-IN PAD

X793 X546-SPLITT-OUT-R-IN X546-SPLITT-OUT-R-INr LSmitll_PTLRX
X794 X546-SPLITT-OUT-R-INr X546-SPLITT-OUT-R-INdc LSmitll_SFQDC
R795 X546-SPLITT-OUT-R-INdc 0 5
X796 X546-SPLITT-OUT-R-IN PAD

X797 X547-SPLITT-OUT-R-IN X547-SPLITT-OUT-R-INr LSmitll_PTLRX
X798 X547-SPLITT-OUT-R-INr X547-SPLITT-OUT-R-INdc LSmitll_SFQDC
R799 X547-SPLITT-OUT-R-INdc 0 5
X800 X547-SPLITT-OUT-R-IN PAD

X801 X548-SPLITT-OUT-R-IN X548-SPLITT-OUT-R-INr LSmitll_PTLRX
X802 X548-SPLITT-OUT-R-INr X548-SPLITT-OUT-R-INdc LSmitll_SFQDC
R803 X548-SPLITT-OUT-R-INdc 0 5
X804 X548-SPLITT-OUT-R-IN PAD

X805 X549-SPLITT-OUT-R-IN X549-SPLITT-OUT-R-INr LSmitll_PTLRX
X806 X549-SPLITT-OUT-R-INr X549-SPLITT-OUT-R-INdc LSmitll_SFQDC
R807 X549-SPLITT-OUT-R-INdc 0 5
X808 X549-SPLITT-OUT-R-IN PAD

X809 X550-SPLITT-OUT-R-IN X550-SPLITT-OUT-R-INr LSmitll_PTLRX
X810 X550-SPLITT-OUT-R-INr X550-SPLITT-OUT-R-INdc LSmitll_SFQDC
R811 X550-SPLITT-OUT-R-INdc 0 5
X812 X550-SPLITT-OUT-R-IN PAD

X813 X551-SPLITT-OUT-R-IN X551-SPLITT-OUT-R-INr LSmitll_PTLRX
X814 X551-SPLITT-OUT-R-INr X551-SPLITT-OUT-R-INdc LSmitll_SFQDC
R815 X551-SPLITT-OUT-R-INdc 0 5
X816 X551-SPLITT-OUT-R-IN PAD

X817 X552-SPLITT-OUT-R-IN X552-SPLITT-OUT-R-INr LSmitll_PTLRX
X818 X552-SPLITT-OUT-R-INr X552-SPLITT-OUT-R-INdc LSmitll_SFQDC
R819 X552-SPLITT-OUT-R-INdc 0 5
X820 X552-SPLITT-OUT-R-IN PAD

X821 X553-SPLITT-OUT-R-IN X553-SPLITT-OUT-R-INr LSmitll_PTLRX
X822 X553-SPLITT-OUT-R-INr X553-SPLITT-OUT-R-INdc LSmitll_SFQDC
R823 X553-SPLITT-OUT-R-INdc 0 5
X824 X553-SPLITT-OUT-R-IN PAD

X825 X554-SPLITT-OUT-R-IN X554-SPLITT-OUT-R-INr LSmitll_PTLRX
X826 X554-SPLITT-OUT-R-INr X554-SPLITT-OUT-R-INdc LSmitll_SFQDC
R827 X554-SPLITT-OUT-R-INdc 0 5
X828 X554-SPLITT-OUT-R-IN PAD

X829 X555-SPLITT-OUT-R-IN X555-SPLITT-OUT-R-INr LSmitll_PTLRX
X830 X555-SPLITT-OUT-R-INr X555-SPLITT-OUT-R-INdc LSmitll_SFQDC
R831 X555-SPLITT-OUT-R-INdc 0 5
X832 X555-SPLITT-OUT-R-IN PAD

X833 X556-SPLITT-OUT-R-IN X556-SPLITT-OUT-R-INr LSmitll_PTLRX
X834 X556-SPLITT-OUT-R-INr X556-SPLITT-OUT-R-INdc LSmitll_SFQDC
R835 X556-SPLITT-OUT-R-INdc 0 5
X836 X556-SPLITT-OUT-R-IN PAD

X837 X557-SPLITT-OUT-R-IN X557-SPLITT-OUT-R-INr LSmitll_PTLRX
X838 X557-SPLITT-OUT-R-INr X557-SPLITT-OUT-R-INdc LSmitll_SFQDC
R839 X557-SPLITT-OUT-R-INdc 0 5
X840 X557-SPLITT-OUT-R-IN PAD

X841 X558-SPLITT-OUT-R-IN X558-SPLITT-OUT-R-INr LSmitll_PTLRX
X842 X558-SPLITT-OUT-R-INr X558-SPLITT-OUT-R-INdc LSmitll_SFQDC
R843 X558-SPLITT-OUT-R-INdc 0 5
X844 X558-SPLITT-OUT-R-IN PAD

X845 X559-SPLITT-OUT-R-IN X559-SPLITT-OUT-R-INr LSmitll_PTLRX
X846 X559-SPLITT-OUT-R-INr X559-SPLITT-OUT-R-INdc LSmitll_SFQDC
R847 X559-SPLITT-OUT-R-INdc 0 5
X848 X559-SPLITT-OUT-R-IN PAD

X849 X560-SPLITT-OUT-R-IN X560-SPLITT-OUT-R-INr LSmitll_PTLRX
X850 X560-SPLITT-OUT-R-INr X560-SPLITT-OUT-R-INdc LSmitll_SFQDC
R851 X560-SPLITT-OUT-R-INdc 0 5
X852 X560-SPLITT-OUT-R-IN PAD

X853 X561-SPLITT-OUT-R-IN X561-SPLITT-OUT-R-INr LSmitll_PTLRX
X854 X561-SPLITT-OUT-R-INr X561-SPLITT-OUT-R-INdc LSmitll_SFQDC
R855 X561-SPLITT-OUT-R-INdc 0 5
X856 X561-SPLITT-OUT-R-IN PAD

X857 X562-SPLITT-OUT-R-IN X562-SPLITT-OUT-R-INr LSmitll_PTLRX
X858 X562-SPLITT-OUT-R-INr X562-SPLITT-OUT-R-INdc LSmitll_SFQDC
R859 X562-SPLITT-OUT-R-INdc 0 5
X860 X562-SPLITT-OUT-R-IN PAD

X861 X563-SPLITT-OUT-R-IN X563-SPLITT-OUT-R-INr LSmitll_PTLRX
X862 X563-SPLITT-OUT-R-INr X563-SPLITT-OUT-R-INdc LSmitll_SFQDC
R863 X563-SPLITT-OUT-R-INdc 0 5
X864 X563-SPLITT-OUT-R-IN PAD



t869 X1-LSmitll_DFFT-OUT-X57-LSmitll_AND2T-INt 0 X1-LSmitll_DFFT-OUT-X57-LSmitll_AND2T-IN 0 z0=5 td=2.9ps
X1 Imm3 X519-LSmitll_SPLITT-OUT-X1-LSmitll_DFFT-IN X1-LSmitll_DFFT-OUT-X57-LSmitll_AND2T-INt LSmitll_DFFT

t870 X2-LSmitll_DFFT-OUT-X59-LSmitll_AND2T-INt 0 X2-LSmitll_DFFT-OUT-X59-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X2 Imm2 X422-LSmitll_SPLITT-OUT-X2-LSmitll_DFFT-IN X2-LSmitll_DFFT-OUT-X59-LSmitll_AND2T-INt LSmitll_DFFT

t871 X3-LSmitll_SPLITT-OUT-X5-LSmitll_SPLITT-INt 0 X3-LSmitll_SPLITT-OUT-X5-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t872 X3-LSmitll_SPLITT-OUT-X4-LSmitll_SPLITT-INt 0 X3-LSmitll_SPLITT-OUT-X4-LSmitll_SPLITT-IN 0 z0=5 td=5.1ps
X3 select1 X3-LSmitll_SPLITT-OUT-X5-LSmitll_SPLITT-INt X3-LSmitll_SPLITT-OUT-X4-LSmitll_SPLITT-INt LSmitll_SPLITT

t873 X4-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-INt 0 X4-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-IN 0 z0=5 td=3.3ps
t874 X4-LSmitll_SPLITT-OUT-X23-LSmitll_NOTT-INt 0 X4-LSmitll_SPLITT-OUT-X23-LSmitll_NOTT-IN 0 z0=5 td=2.2ps
X4 X3-LSmitll_SPLITT-OUT-X4-LSmitll_SPLITT-IN X4-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-INt X4-LSmitll_SPLITT-OUT-X23-LSmitll_NOTT-INt LSmitll_SPLITT

t875 X5-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-INt 0 X5-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
t876 X5-LSmitll_SPLITT-OUT-X25-LSmitll_NOTT-INt 0 X5-LSmitll_SPLITT-OUT-X25-LSmitll_NOTT-IN 0 z0=5 td=1.1ps
X5 X3-LSmitll_SPLITT-OUT-X5-LSmitll_SPLITT-IN X5-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-INt X5-LSmitll_SPLITT-OUT-X25-LSmitll_NOTT-INt LSmitll_SPLITT

t877 X6-LSmitll_DFFT-OUT-X61-LSmitll_AND2T-INt 0 X6-LSmitll_DFFT-OUT-X61-LSmitll_AND2T-IN 0 z0=5 td=11.3ps
X6 Imm1 X342-LSmitll_SPLITT-OUT-X6-LSmitll_DFFT-IN X6-LSmitll_DFFT-OUT-X61-LSmitll_AND2T-INt LSmitll_DFFT

t878 X7-LSmitll_DFFT-OUT-X63-LSmitll_AND2T-INt 0 X7-LSmitll_DFFT-OUT-X63-LSmitll_AND2T-IN 0 z0=5 td=2.7ps
X7 Imm0 X520-LSmitll_SPLITT-OUT-X7-LSmitll_DFFT-IN X7-LSmitll_DFFT-OUT-X63-LSmitll_AND2T-INt LSmitll_DFFT

t879 X8-LSmitll_SPLITT-OUT-X10-LSmitll_SPLITT-INt 0 X8-LSmitll_SPLITT-OUT-X10-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t880 X8-LSmitll_SPLITT-OUT-X9-LSmitll_SPLITT-INt 0 X8-LSmitll_SPLITT-OUT-X9-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X8 select0 X8-LSmitll_SPLITT-OUT-X10-LSmitll_SPLITT-INt X8-LSmitll_SPLITT-OUT-X9-LSmitll_SPLITT-INt LSmitll_SPLITT

t881 X9-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-INt 0 X9-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-IN 0 z0=5 td=3.2ps
t882 X9-LSmitll_SPLITT-OUT-X27-LSmitll_NOTT-INt 0 X9-LSmitll_SPLITT-OUT-X27-LSmitll_NOTT-IN 0 z0=5 td=1.1ps
X9 X8-LSmitll_SPLITT-OUT-X9-LSmitll_SPLITT-IN X9-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-INt X9-LSmitll_SPLITT-OUT-X27-LSmitll_NOTT-INt LSmitll_SPLITT

t883 X10-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-INt 0 X10-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t884 X10-LSmitll_SPLITT-OUT-X29-LSmitll_NOTT-INt 0 X10-LSmitll_SPLITT-OUT-X29-LSmitll_NOTT-IN 0 z0=5 td=10.9ps
X10 X8-LSmitll_SPLITT-OUT-X10-LSmitll_SPLITT-IN X10-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-INt X10-LSmitll_SPLITT-OUT-X29-LSmitll_NOTT-INt LSmitll_SPLITT

t885 X11-LSmitll_SPLITT-OUT-X13-LSmitll_SPLITT-INt 0 X11-LSmitll_SPLITT-OUT-X13-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t886 X11-LSmitll_SPLITT-OUT-X12-LSmitll_SPLITT-INt 0 X11-LSmitll_SPLITT-OUT-X12-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X11 read X11-LSmitll_SPLITT-OUT-X13-LSmitll_SPLITT-INt X11-LSmitll_SPLITT-OUT-X12-LSmitll_SPLITT-INt LSmitll_SPLITT

t887 X12-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-INt 0 X12-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-IN 0 z0=5 td=3.1ps
t888 X12-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-INt 0 X12-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
X12 X11-LSmitll_SPLITT-OUT-X12-LSmitll_SPLITT-IN X12-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-INt X12-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-INt LSmitll_SPLITT

t889 X13-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-INt 0 X13-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-IN 0 z0=5 td=3.3ps
t890 X13-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-INt 0 X13-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X13 X11-LSmitll_SPLITT-OUT-X13-LSmitll_SPLITT-IN X13-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-INt X13-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-INt LSmitll_SPLITT

t891 X14-LSmitll_SPLITT-OUT-X36-LSmitll_DFFT-INt 0 X14-LSmitll_SPLITT-OUT-X36-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
t892 X14-LSmitll_SPLITT-OUT-X35-LSmitll_DFFT-INt 0 X14-LSmitll_SPLITT-OUT-X35-LSmitll_DFFT-IN 0 z0=5 td=3.9ps
X14 addr0 X14-LSmitll_SPLITT-OUT-X36-LSmitll_DFFT-INt X14-LSmitll_SPLITT-OUT-X35-LSmitll_DFFT-INt LSmitll_SPLITT

t893 X15-LSmitll_SPLITT-OUT-X38-LSmitll_DFFT-INt 0 X15-LSmitll_SPLITT-OUT-X38-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t894 X15-LSmitll_SPLITT-OUT-X37-LSmitll_DFFT-INt 0 X15-LSmitll_SPLITT-OUT-X37-LSmitll_DFFT-IN 0 z0=5 td=2.7ps
X15 addr1 X15-LSmitll_SPLITT-OUT-X38-LSmitll_DFFT-INt X15-LSmitll_SPLITT-OUT-X37-LSmitll_DFFT-INt LSmitll_SPLITT

t895 X16-LSmitll_SPLITT-OUT-X40-LSmitll_DFFT-INt 0 X16-LSmitll_SPLITT-OUT-X40-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t896 X16-LSmitll_SPLITT-OUT-X39-LSmitll_DFFT-INt 0 X16-LSmitll_SPLITT-OUT-X39-LSmitll_DFFT-IN 0 z0=5 td=4.5ps
X16 write_flags X16-LSmitll_SPLITT-OUT-X40-LSmitll_DFFT-INt X16-LSmitll_SPLITT-OUT-X39-LSmitll_DFFT-INt LSmitll_SPLITT

t897 X17-LSmitll_SPLITT-OUT-X143-LSmitll_XORT-INt 0 X17-LSmitll_SPLITT-OUT-X143-LSmitll_XORT-IN 0 z0=5 td=2.1ps
t898 X17-LSmitll_SPLITT-OUT-X141-LSmitll_XORT-INt 0 X17-LSmitll_SPLITT-OUT-X141-LSmitll_XORT-IN 0 z0=5 td=2.7ps
X17 Cmpl_b1 X17-LSmitll_SPLITT-OUT-X143-LSmitll_XORT-INt X17-LSmitll_SPLITT-OUT-X141-LSmitll_XORT-INt LSmitll_SPLITT

t899 X18-LSmitll_SPLITT-OUT-X147-LSmitll_XORT-INt 0 X18-LSmitll_SPLITT-OUT-X147-LSmitll_XORT-IN 0 z0=5 td=3.2ps
t900 X18-LSmitll_SPLITT-OUT-X145-LSmitll_XORT-INt 0 X18-LSmitll_SPLITT-OUT-X145-LSmitll_XORT-IN 0 z0=5 td=2.2ps
X18 Cmpl_b0 X18-LSmitll_SPLITT-OUT-X147-LSmitll_XORT-INt X18-LSmitll_SPLITT-OUT-X145-LSmitll_XORT-INt LSmitll_SPLITT

t901 X19-LSmitll_DFFT-OUT-X167-LSmitll_DFFT-INt 0 X19-LSmitll_DFFT-OUT-X167-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X19 Cin X362-LSmitll_SPLITT-OUT-X19-LSmitll_DFFT-IN X19-LSmitll_DFFT-OUT-X167-LSmitll_DFFT-INt LSmitll_DFFT

t902 X20-LSmitll_DFFT-OUT-X164-LSmitll_DFFT-INt 0 X20-LSmitll_DFFT-OUT-X164-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X20 Op_Arith X323-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-IN X20-LSmitll_DFFT-OUT-X164-LSmitll_DFFT-INt LSmitll_DFFT

t903 X21-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-INt 0 X21-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X21 Op_And X521-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-IN X21-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-INt LSmitll_DFFT

t904 X22-LSmitll_DFFT-OUT-X166-LSmitll_DFFT-INt 0 X22-LSmitll_DFFT-OUT-X166-LSmitll_DFFT-IN 0 z0=5 td=3.5ps
X22 Op_Xor X375-LSmitll_SPLITT-OUT-X22-LSmitll_DFFT-IN X22-LSmitll_DFFT-OUT-X166-LSmitll_DFFT-INt LSmitll_DFFT

t905 X23-LSmitll_NOTT-OUT-X57-LSmitll_AND2T-INt 0 X23-LSmitll_NOTT-OUT-X57-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
X23 X4-LSmitll_SPLITT-OUT-X23-LSmitll_NOTT-IN X441-LSmitll_SPLITT-OUT-X23-LSmitll_NOTT-IN X23-LSmitll_NOTT-OUT-X57-LSmitll_AND2T-INt LSmitll_NOTT

t906 X24-LSmitll_DFFT-OUT-X58-LSmitll_AND2T-INt 0 X24-LSmitll_DFFT-OUT-X58-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
X24 X4-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-IN X441-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-IN X24-LSmitll_DFFT-OUT-X58-LSmitll_AND2T-INt LSmitll_DFFT

t907 X25-LSmitll_NOTT-OUT-X59-LSmitll_AND2T-INt 0 X25-LSmitll_NOTT-OUT-X59-LSmitll_AND2T-IN 0 z0=5 td=4.7ps
X25 X5-LSmitll_SPLITT-OUT-X25-LSmitll_NOTT-IN X415-LSmitll_SPLITT-OUT-X25-LSmitll_NOTT-IN X25-LSmitll_NOTT-OUT-X59-LSmitll_AND2T-INt LSmitll_NOTT

t908 X26-LSmitll_DFFT-OUT-X60-LSmitll_AND2T-INt 0 X26-LSmitll_DFFT-OUT-X60-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
X26 X5-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-IN X421-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-IN X26-LSmitll_DFFT-OUT-X60-LSmitll_AND2T-INt LSmitll_DFFT

t909 X27-LSmitll_NOTT-OUT-X61-LSmitll_AND2T-INt 0 X27-LSmitll_NOTT-OUT-X61-LSmitll_AND2T-IN 0 z0=5 td=14.8ps
X27 X9-LSmitll_SPLITT-OUT-X27-LSmitll_NOTT-IN X317-LSmitll_SPLITT-OUT-X27-LSmitll_NOTT-IN X27-LSmitll_NOTT-OUT-X61-LSmitll_AND2T-INt LSmitll_NOTT

t910 X28-LSmitll_DFFT-OUT-X62-LSmitll_AND2T-INt 0 X28-LSmitll_DFFT-OUT-X62-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X28 X9-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-IN X311-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-IN X28-LSmitll_DFFT-OUT-X62-LSmitll_AND2T-INt LSmitll_DFFT

t911 X29-LSmitll_NOTT-OUT-X63-LSmitll_AND2T-INt 0 X29-LSmitll_NOTT-OUT-X63-LSmitll_AND2T-IN 0 z0=5 td=3.8ps
X29 X10-LSmitll_SPLITT-OUT-X29-LSmitll_NOTT-IN X337-LSmitll_SPLITT-OUT-X29-LSmitll_NOTT-IN X29-LSmitll_NOTT-OUT-X63-LSmitll_AND2T-INt LSmitll_NOTT

t912 X30-LSmitll_DFFT-OUT-X64-LSmitll_AND2T-INt 0 X30-LSmitll_DFFT-OUT-X64-LSmitll_AND2T-IN 0 z0=5 td=12.1ps
X30 X10-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-IN X336-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-IN X30-LSmitll_DFFT-OUT-X64-LSmitll_AND2T-INt LSmitll_DFFT

t913 X31-LSmitll_DFFT-OUT-X65-LSmitll_DFFT-INt 0 X31-LSmitll_DFFT-OUT-X65-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X31 X12-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-IN X403-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-IN X31-LSmitll_DFFT-OUT-X65-LSmitll_DFFT-INt LSmitll_DFFT

t914 X32-LSmitll_DFFT-OUT-X66-LSmitll_DFFT-INt 0 X32-LSmitll_DFFT-OUT-X66-LSmitll_DFFT-IN 0 z0=5 td=14.8ps
X32 X12-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-IN X408-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-IN X32-LSmitll_DFFT-OUT-X66-LSmitll_DFFT-INt LSmitll_DFFT

t915 X33-LSmitll_DFFT-OUT-X67-LSmitll_DFFT-INt 0 X33-LSmitll_DFFT-OUT-X67-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X33 X13-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-IN X406-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-IN X33-LSmitll_DFFT-OUT-X67-LSmitll_DFFT-INt LSmitll_DFFT

t916 X34-LSmitll_DFFT-OUT-X68-LSmitll_DFFT-INt 0 X34-LSmitll_DFFT-OUT-X68-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X34 X13-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-IN X522-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-IN X34-LSmitll_DFFT-OUT-X68-LSmitll_DFFT-INt LSmitll_DFFT

t917 X35-LSmitll_DFFT-OUT-X41-LSmitll_SPLITT-INt 0 X35-LSmitll_DFFT-OUT-X41-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X35 X14-LSmitll_SPLITT-OUT-X35-LSmitll_DFFT-IN X344-LSmitll_SPLITT-OUT-X35-LSmitll_DFFT-IN X35-LSmitll_DFFT-OUT-X41-LSmitll_SPLITT-INt LSmitll_DFFT

t918 X36-LSmitll_DFFT-OUT-X44-LSmitll_SPLITT-INt 0 X36-LSmitll_DFFT-OUT-X44-LSmitll_SPLITT-IN 0 z0=5 td=11.6ps
X36 X14-LSmitll_SPLITT-OUT-X36-LSmitll_DFFT-IN X317-LSmitll_SPLITT-OUT-X36-LSmitll_DFFT-IN X36-LSmitll_DFFT-OUT-X44-LSmitll_SPLITT-INt LSmitll_DFFT

t919 X37-LSmitll_DFFT-OUT-X47-LSmitll_SPLITT-INt 0 X37-LSmitll_DFFT-OUT-X47-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X37 X15-LSmitll_SPLITT-OUT-X37-LSmitll_DFFT-IN X313-LSmitll_SPLITT-OUT-X37-LSmitll_DFFT-IN X37-LSmitll_DFFT-OUT-X47-LSmitll_SPLITT-INt LSmitll_DFFT

t920 X38-LSmitll_DFFT-OUT-X50-LSmitll_SPLITT-INt 0 X38-LSmitll_DFFT-OUT-X50-LSmitll_SPLITT-IN 0 z0=5 td=4.8ps
X38 X15-LSmitll_SPLITT-OUT-X38-LSmitll_DFFT-IN X313-LSmitll_SPLITT-OUT-X38-LSmitll_DFFT-IN X38-LSmitll_DFFT-OUT-X50-LSmitll_SPLITT-INt LSmitll_DFFT

t921 X39-LSmitll_DFFT-OUT-X54-LSmitll_SPLITT-INt 0 X39-LSmitll_DFFT-OUT-X54-LSmitll_SPLITT-IN 0 z0=5 td=8.9ps
X39 X16-LSmitll_SPLITT-OUT-X39-LSmitll_DFFT-IN X444-LSmitll_SPLITT-OUT-X39-LSmitll_DFFT-IN X39-LSmitll_DFFT-OUT-X54-LSmitll_SPLITT-INt LSmitll_DFFT

t922 X40-LSmitll_DFFT-OUT-X53-LSmitll_SPLITT-INt 0 X40-LSmitll_DFFT-OUT-X53-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X40 X16-LSmitll_SPLITT-OUT-X40-LSmitll_DFFT-IN X344-LSmitll_SPLITT-OUT-X40-LSmitll_DFFT-IN X40-LSmitll_DFFT-OUT-X53-LSmitll_SPLITT-INt LSmitll_DFFT

t923 X41-LSmitll_SPLITT-OUT-X43-LSmitll_SPLITT-INt 0 X41-LSmitll_SPLITT-OUT-X43-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t924 X41-LSmitll_SPLITT-OUT-X42-LSmitll_SPLITT-INt 0 X41-LSmitll_SPLITT-OUT-X42-LSmitll_SPLITT-IN 0 z0=5 td=3.5ps
X41 X35-LSmitll_DFFT-OUT-X41-LSmitll_SPLITT-IN X41-LSmitll_SPLITT-OUT-X43-LSmitll_SPLITT-INt X41-LSmitll_SPLITT-OUT-X42-LSmitll_SPLITT-INt LSmitll_SPLITT

t925 X42-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-INt 0 X42-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
t926 X42-LSmitll_SPLITT-OUT-X85-LSmitll_NDROT-INt 0 X42-LSmitll_SPLITT-OUT-X85-LSmitll_NDROT-IN 0 z0=5 td=2.4ps
X42 X41-LSmitll_SPLITT-OUT-X42-LSmitll_SPLITT-IN X42-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-INt X42-LSmitll_SPLITT-OUT-X85-LSmitll_NDROT-INt LSmitll_SPLITT

t927 X43-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-INt 0 X43-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t928 X43-LSmitll_SPLITT-OUT-X88-LSmitll_NDROT-INt 0 X43-LSmitll_SPLITT-OUT-X88-LSmitll_NDROT-IN 0 z0=5 td=2.8ps
X43 X41-LSmitll_SPLITT-OUT-X43-LSmitll_SPLITT-IN X43-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-INt X43-LSmitll_SPLITT-OUT-X88-LSmitll_NDROT-INt LSmitll_SPLITT

t929 X44-LSmitll_SPLITT-OUT-X46-LSmitll_SPLITT-INt 0 X44-LSmitll_SPLITT-OUT-X46-LSmitll_SPLITT-IN 0 z0=5 td=3.2ps
t930 X44-LSmitll_SPLITT-OUT-X45-LSmitll_SPLITT-INt 0 X44-LSmitll_SPLITT-OUT-X45-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X44 X36-LSmitll_DFFT-OUT-X44-LSmitll_SPLITT-IN X44-LSmitll_SPLITT-OUT-X46-LSmitll_SPLITT-INt X44-LSmitll_SPLITT-OUT-X45-LSmitll_SPLITT-INt LSmitll_SPLITT

t931 X45-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-INt 0 X45-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-IN 0 z0=5 td=4.5ps
t932 X45-LSmitll_SPLITT-OUT-X91-LSmitll_NDROT-INt 0 X45-LSmitll_SPLITT-OUT-X91-LSmitll_NDROT-IN 0 z0=5 td=1.1ps
X45 X44-LSmitll_SPLITT-OUT-X45-LSmitll_SPLITT-IN X45-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-INt X45-LSmitll_SPLITT-OUT-X91-LSmitll_NDROT-INt LSmitll_SPLITT

t933 X46-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-INt 0 X46-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-IN 0 z0=5 td=2.7ps
t934 X46-LSmitll_SPLITT-OUT-X94-LSmitll_NDROT-INt 0 X46-LSmitll_SPLITT-OUT-X94-LSmitll_NDROT-IN 0 z0=5 td=5.7ps
X46 X44-LSmitll_SPLITT-OUT-X46-LSmitll_SPLITT-IN X46-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-INt X46-LSmitll_SPLITT-OUT-X94-LSmitll_NDROT-INt LSmitll_SPLITT

t935 X47-LSmitll_SPLITT-OUT-X49-LSmitll_SPLITT-INt 0 X47-LSmitll_SPLITT-OUT-X49-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t936 X47-LSmitll_SPLITT-OUT-X48-LSmitll_SPLITT-INt 0 X47-LSmitll_SPLITT-OUT-X48-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X47 X37-LSmitll_DFFT-OUT-X47-LSmitll_SPLITT-IN X47-LSmitll_SPLITT-OUT-X49-LSmitll_SPLITT-INt X47-LSmitll_SPLITT-OUT-X48-LSmitll_SPLITT-INt LSmitll_SPLITT

t937 X48-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-INt 0 X48-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-IN 0 z0=5 td=3.4ps
t938 X48-LSmitll_SPLITT-OUT-X97-LSmitll_NDROT-INt 0 X48-LSmitll_SPLITT-OUT-X97-LSmitll_NDROT-IN 0 z0=5 td=2.4ps
X48 X47-LSmitll_SPLITT-OUT-X48-LSmitll_SPLITT-IN X48-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-INt X48-LSmitll_SPLITT-OUT-X97-LSmitll_NDROT-INt LSmitll_SPLITT

t939 X49-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt 0 X49-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t940 X49-LSmitll_SPLITT-OUT-X100-LSmitll_NDROT-INt 0 X49-LSmitll_SPLITT-OUT-X100-LSmitll_NDROT-IN 0 z0=5 td=1.1ps
X49 X47-LSmitll_SPLITT-OUT-X49-LSmitll_SPLITT-IN X49-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt X49-LSmitll_SPLITT-OUT-X100-LSmitll_NDROT-INt LSmitll_SPLITT

t941 X50-LSmitll_SPLITT-OUT-X52-LSmitll_SPLITT-INt 0 X50-LSmitll_SPLITT-OUT-X52-LSmitll_SPLITT-IN 0 z0=5 td=3.7ps
t942 X50-LSmitll_SPLITT-OUT-X51-LSmitll_SPLITT-INt 0 X50-LSmitll_SPLITT-OUT-X51-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X50 X38-LSmitll_DFFT-OUT-X50-LSmitll_SPLITT-IN X50-LSmitll_SPLITT-OUT-X52-LSmitll_SPLITT-INt X50-LSmitll_SPLITT-OUT-X51-LSmitll_SPLITT-INt LSmitll_SPLITT

t943 X51-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt 0 X51-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN 0 z0=5 td=3.6ps
t944 X51-LSmitll_SPLITT-OUT-X103-LSmitll_NDROT-INt 0 X51-LSmitll_SPLITT-OUT-X103-LSmitll_NDROT-IN 0 z0=5 td=2.4ps
X51 X50-LSmitll_SPLITT-OUT-X51-LSmitll_SPLITT-IN X51-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt X51-LSmitll_SPLITT-OUT-X103-LSmitll_NDROT-INt LSmitll_SPLITT

t945 X52-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt 0 X52-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t946 X52-LSmitll_SPLITT-OUT-X106-LSmitll_NDROT-INt 0 X52-LSmitll_SPLITT-OUT-X106-LSmitll_NDROT-IN 0 z0=5 td=4.1ps
X52 X50-LSmitll_SPLITT-OUT-X52-LSmitll_SPLITT-IN X52-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt X52-LSmitll_SPLITT-OUT-X106-LSmitll_NDROT-INt LSmitll_SPLITT

t947 X53-LSmitll_SPLITT-OUT-X116-LSmitll_AND2T-INt 0 X53-LSmitll_SPLITT-OUT-X116-LSmitll_AND2T-IN 0 z0=5 td=3.6ps
t948 X53-LSmitll_SPLITT-OUT-X115-LSmitll_NDROT-INt 0 X53-LSmitll_SPLITT-OUT-X115-LSmitll_NDROT-IN 0 z0=5 td=2.4ps
X53 X40-LSmitll_DFFT-OUT-X53-LSmitll_SPLITT-IN X53-LSmitll_SPLITT-OUT-X116-LSmitll_AND2T-INt X53-LSmitll_SPLITT-OUT-X115-LSmitll_NDROT-INt LSmitll_SPLITT

t949 X54-LSmitll_SPLITT-OUT-X56-LSmitll_SPLITT-INt 0 X54-LSmitll_SPLITT-OUT-X56-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t950 X54-LSmitll_SPLITT-OUT-X55-LSmitll_SPLITT-INt 0 X54-LSmitll_SPLITT-OUT-X55-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X54 X39-LSmitll_DFFT-OUT-X54-LSmitll_SPLITT-IN X54-LSmitll_SPLITT-OUT-X56-LSmitll_SPLITT-INt X54-LSmitll_SPLITT-OUT-X55-LSmitll_SPLITT-INt LSmitll_SPLITT

t951 X55-LSmitll_SPLITT-OUT-X110-LSmitll_AND2T-INt 0 X55-LSmitll_SPLITT-OUT-X110-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t952 X55-LSmitll_SPLITT-OUT-X109-LSmitll_NDROT-INt 0 X55-LSmitll_SPLITT-OUT-X109-LSmitll_NDROT-IN 0 z0=5 td=7.7ps
X55 X54-LSmitll_SPLITT-OUT-X55-LSmitll_SPLITT-IN X55-LSmitll_SPLITT-OUT-X110-LSmitll_AND2T-INt X55-LSmitll_SPLITT-OUT-X109-LSmitll_NDROT-INt LSmitll_SPLITT

t953 X56-LSmitll_SPLITT-OUT-X113-LSmitll_AND2T-INt 0 X56-LSmitll_SPLITT-OUT-X113-LSmitll_AND2T-IN 0 z0=5 td=4.2ps
t954 X56-LSmitll_SPLITT-OUT-X112-LSmitll_NDROT-INt 0 X56-LSmitll_SPLITT-OUT-X112-LSmitll_NDROT-IN 0 z0=5 td=2.4ps
X56 X54-LSmitll_SPLITT-OUT-X56-LSmitll_SPLITT-IN X56-LSmitll_SPLITT-OUT-X113-LSmitll_AND2T-INt X56-LSmitll_SPLITT-OUT-X112-LSmitll_NDROT-INt LSmitll_SPLITT

t955 X57-LSmitll_AND2T-OUT-X73-LSmitll_OR2T-INt 0 X57-LSmitll_AND2T-OUT-X73-LSmitll_OR2T-IN 0 z0=5 td=2.6ps
X57 X1-LSmitll_DFFT-OUT-X57-LSmitll_AND2T-IN X23-LSmitll_NOTT-OUT-X57-LSmitll_AND2T-IN X442-LSmitll_SPLITT-OUT-X57-LSmitll_AND2T-IN X57-LSmitll_AND2T-OUT-X73-LSmitll_OR2T-INt LSmitll_AND2T

t956 X58-LSmitll_AND2T-OUT-X73-LSmitll_OR2T-INt 0 X58-LSmitll_AND2T-OUT-X73-LSmitll_OR2T-IN 0 z0=5 td=4.3ps
X58 X24-LSmitll_DFFT-OUT-X58-LSmitll_AND2T-IN X303-LSmitll_DFFT-OUT-X58-LSmitll_AND2T-IN X442-LSmitll_SPLITT-OUT-X58-LSmitll_AND2T-IN X58-LSmitll_AND2T-OUT-X73-LSmitll_OR2T-INt LSmitll_AND2T

t957 X59-LSmitll_AND2T-OUT-X74-LSmitll_OR2T-INt 0 X59-LSmitll_AND2T-OUT-X74-LSmitll_OR2T-IN 0 z0=5 td=2.4ps
X59 X2-LSmitll_DFFT-OUT-X59-LSmitll_AND2T-IN X25-LSmitll_NOTT-OUT-X59-LSmitll_AND2T-IN X421-LSmitll_SPLITT-OUT-X59-LSmitll_AND2T-IN X59-LSmitll_AND2T-OUT-X74-LSmitll_OR2T-INt LSmitll_AND2T

t958 X60-LSmitll_AND2T-OUT-X74-LSmitll_OR2T-INt 0 X60-LSmitll_AND2T-OUT-X74-LSmitll_OR2T-IN 0 z0=5 td=2.9ps
X60 X26-LSmitll_DFFT-OUT-X60-LSmitll_AND2T-IN X304-LSmitll_DFFT-OUT-X60-LSmitll_AND2T-IN X422-LSmitll_SPLITT-OUT-X60-LSmitll_AND2T-IN X60-LSmitll_AND2T-OUT-X74-LSmitll_OR2T-INt LSmitll_AND2T

t959 X61-LSmitll_AND2T-OUT-X75-LSmitll_OR2T-INt 0 X61-LSmitll_AND2T-OUT-X75-LSmitll_OR2T-IN 0 z0=5 td=2.6ps
X61 X6-LSmitll_DFFT-OUT-X61-LSmitll_AND2T-IN X27-LSmitll_NOTT-OUT-X61-LSmitll_AND2T-IN X310-LSmitll_SPLITT-OUT-X61-LSmitll_AND2T-IN X61-LSmitll_AND2T-OUT-X75-LSmitll_OR2T-INt LSmitll_AND2T

t960 X62-LSmitll_AND2T-OUT-X75-LSmitll_OR2T-INt 0 X62-LSmitll_AND2T-OUT-X75-LSmitll_OR2T-IN 0 z0=5 td=1.4ps
X62 X28-LSmitll_DFFT-OUT-X62-LSmitll_AND2T-IN X305-LSmitll_DFFT-OUT-X62-LSmitll_AND2T-IN X311-LSmitll_SPLITT-OUT-X62-LSmitll_AND2T-IN X62-LSmitll_AND2T-OUT-X75-LSmitll_OR2T-INt LSmitll_AND2T

t961 X63-LSmitll_AND2T-OUT-X76-LSmitll_OR2T-INt 0 X63-LSmitll_AND2T-OUT-X76-LSmitll_OR2T-IN 0 z0=5 td=2.6ps
X63 X7-LSmitll_DFFT-OUT-X63-LSmitll_AND2T-IN X29-LSmitll_NOTT-OUT-X63-LSmitll_AND2T-IN X523-LSmitll_SPLITT-OUT-X63-LSmitll_AND2T-IN X63-LSmitll_AND2T-OUT-X76-LSmitll_OR2T-INt LSmitll_AND2T

t962 X64-LSmitll_AND2T-OUT-X76-LSmitll_OR2T-INt 0 X64-LSmitll_AND2T-OUT-X76-LSmitll_OR2T-IN 0 z0=5 td=4.5ps
X64 X30-LSmitll_DFFT-OUT-X64-LSmitll_AND2T-IN X306-LSmitll_DFFT-OUT-X64-LSmitll_AND2T-IN X342-LSmitll_SPLITT-OUT-X64-LSmitll_AND2T-IN X64-LSmitll_AND2T-OUT-X76-LSmitll_OR2T-INt LSmitll_AND2T

t963 X65-LSmitll_DFFT-OUT-X69-LSmitll_SPLITT-INt 0 X65-LSmitll_DFFT-OUT-X69-LSmitll_SPLITT-IN 0 z0=5 td=11.7ps
X65 X31-LSmitll_DFFT-OUT-X65-LSmitll_DFFT-IN X524-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-IN X65-LSmitll_DFFT-OUT-X69-LSmitll_SPLITT-INt LSmitll_DFFT

t964 X66-LSmitll_DFFT-OUT-X70-LSmitll_SPLITT-INt 0 X66-LSmitll_DFFT-OUT-X70-LSmitll_SPLITT-IN 0 z0=5 td=4.7ps
X66 X32-LSmitll_DFFT-OUT-X66-LSmitll_DFFT-IN X507-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-IN X66-LSmitll_DFFT-OUT-X70-LSmitll_SPLITT-INt LSmitll_DFFT

t965 X67-LSmitll_DFFT-OUT-X71-LSmitll_SPLITT-INt 0 X67-LSmitll_DFFT-OUT-X71-LSmitll_SPLITT-IN 0 z0=5 td=7.2ps
X67 X33-LSmitll_DFFT-OUT-X67-LSmitll_DFFT-IN X525-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-IN X67-LSmitll_DFFT-OUT-X71-LSmitll_SPLITT-INt LSmitll_DFFT

t966 X68-LSmitll_DFFT-OUT-X72-LSmitll_SPLITT-INt 0 X68-LSmitll_DFFT-OUT-X72-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X68 X34-LSmitll_DFFT-OUT-X68-LSmitll_DFFT-IN X487-LSmitll_SPLITT-OUT-X68-LSmitll_DFFT-IN X68-LSmitll_DFFT-OUT-X72-LSmitll_SPLITT-INt LSmitll_DFFT

t967 X69-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt 0 X69-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN 0 z0=5 td=3.3ps
t968 X69-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-INt 0 X69-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-IN 0 z0=5 td=3.6ps
X69 X65-LSmitll_DFFT-OUT-X69-LSmitll_SPLITT-IN X69-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt X69-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-INt LSmitll_SPLITT

t969 X70-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt 0 X70-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN 0 z0=5 td=3.7ps
t970 X70-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt 0 X70-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN 0 z0=5 td=3.9ps
X70 X66-LSmitll_DFFT-OUT-X70-LSmitll_SPLITT-IN X70-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt X70-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt LSmitll_SPLITT

t971 X71-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-INt 0 X71-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-IN 0 z0=5 td=4.1ps
t972 X71-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt 0 X71-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN 0 z0=5 td=1.9ps
X71 X67-LSmitll_DFFT-OUT-X71-LSmitll_SPLITT-IN X71-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-INt X71-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt LSmitll_SPLITT

t973 X72-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt 0 X72-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN 0 z0=5 td=6.0ps
t974 X72-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt 0 X72-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN 0 z0=5 td=3.0ps
X72 X68-LSmitll_DFFT-OUT-X72-LSmitll_SPLITT-IN X72-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt X72-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt LSmitll_SPLITT

t975 X73-LSmitll_OR2T-OUT-X78-LSmitll_DFFT-INt 0 X73-LSmitll_OR2T-OUT-X78-LSmitll_DFFT-IN 0 z0=5 td=5.2ps
X73 X57-LSmitll_AND2T-OUT-X73-LSmitll_OR2T-IN X58-LSmitll_AND2T-OUT-X73-LSmitll_OR2T-IN X447-LSmitll_SPLITT-OUT-X73-LSmitll_OR2T-IN X73-LSmitll_OR2T-OUT-X78-LSmitll_DFFT-INt LSmitll_OR2T

t976 X74-LSmitll_OR2T-OUT-X77-LSmitll_DFFT-INt 0 X74-LSmitll_OR2T-OUT-X77-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X74 X59-LSmitll_AND2T-OUT-X74-LSmitll_OR2T-IN X60-LSmitll_AND2T-OUT-X74-LSmitll_OR2T-IN X416-LSmitll_SPLITT-OUT-X74-LSmitll_OR2T-IN X74-LSmitll_OR2T-OUT-X77-LSmitll_DFFT-INt LSmitll_OR2T

t977 X75-LSmitll_OR2T-OUT-X80-LSmitll_DFFT-INt 0 X75-LSmitll_OR2T-OUT-X80-LSmitll_DFFT-IN 0 z0=5 td=4.2ps
X75 X61-LSmitll_AND2T-OUT-X75-LSmitll_OR2T-IN X62-LSmitll_AND2T-OUT-X75-LSmitll_OR2T-IN X310-LSmitll_SPLITT-OUT-X75-LSmitll_OR2T-IN X75-LSmitll_OR2T-OUT-X80-LSmitll_DFFT-INt LSmitll_OR2T

t978 X76-LSmitll_OR2T-OUT-X79-LSmitll_DFFT-INt 0 X76-LSmitll_OR2T-OUT-X79-LSmitll_DFFT-IN 0 z0=5 td=6.0ps
X76 X63-LSmitll_AND2T-OUT-X76-LSmitll_OR2T-IN X64-LSmitll_AND2T-OUT-X76-LSmitll_OR2T-IN X415-LSmitll_SPLITT-OUT-X76-LSmitll_OR2T-IN X76-LSmitll_OR2T-OUT-X79-LSmitll_DFFT-INt LSmitll_OR2T

t979 X77-LSmitll_DFFT-OUT-X81-LSmitll_SPLITT-INt 0 X77-LSmitll_DFFT-OUT-X81-LSmitll_SPLITT-IN 0 z0=5 td=5.0ps
X77 X74-LSmitll_OR2T-OUT-X77-LSmitll_DFFT-IN X416-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-IN X77-LSmitll_DFFT-OUT-X81-LSmitll_SPLITT-INt LSmitll_DFFT

t980 X78-LSmitll_DFFT-OUT-X82-LSmitll_SPLITT-INt 0 X78-LSmitll_DFFT-OUT-X82-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X78 X73-LSmitll_OR2T-OUT-X78-LSmitll_DFFT-IN X444-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-IN X78-LSmitll_DFFT-OUT-X82-LSmitll_SPLITT-INt LSmitll_DFFT

t981 X79-LSmitll_DFFT-OUT-X83-LSmitll_SPLITT-INt 0 X79-LSmitll_DFFT-OUT-X83-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
X79 X76-LSmitll_OR2T-OUT-X79-LSmitll_DFFT-IN X339-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-IN X79-LSmitll_DFFT-OUT-X83-LSmitll_SPLITT-INt LSmitll_DFFT

t982 X80-LSmitll_DFFT-OUT-X84-LSmitll_SPLITT-INt 0 X80-LSmitll_DFFT-OUT-X84-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X80 X75-LSmitll_OR2T-OUT-X80-LSmitll_DFFT-IN X526-LSmitll_SPLITT-OUT-X80-LSmitll_DFFT-IN X80-LSmitll_DFFT-OUT-X84-LSmitll_SPLITT-INt LSmitll_DFFT

t983 X81-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt 0 X81-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN 0 z0=5 td=2.6ps
t984 X81-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-INt 0 X81-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X81 X77-LSmitll_DFFT-OUT-X81-LSmitll_SPLITT-IN X81-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt X81-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-INt LSmitll_SPLITT

t985 X82-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt 0 X82-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t986 X82-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-INt 0 X82-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X82 X78-LSmitll_DFFT-OUT-X82-LSmitll_SPLITT-IN X82-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt X82-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-INt LSmitll_SPLITT

t987 X83-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-INt 0 X83-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-IN 0 z0=5 td=3.9ps
t988 X83-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-INt 0 X83-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-IN 0 z0=5 td=5.6ps
X83 X79-LSmitll_DFFT-OUT-X83-LSmitll_SPLITT-IN X83-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-INt X83-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-INt LSmitll_SPLITT

t989 X84-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt 0 X84-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
t990 X84-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-INt 0 X84-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-IN 0 z0=5 td=4.0ps
X84 X80-LSmitll_DFFT-OUT-X84-LSmitll_SPLITT-IN X84-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt X84-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-INt LSmitll_SPLITT

t991 X85-LSmitll_NDROT-OUT-X87-LSmitll_SPLITT-INt 0 X85-LSmitll_NDROT-OUT-X87-LSmitll_SPLITT-IN 0 z0=5 td=6.3ps
X85 X86-LSmitll_AND2T-OUT-X85-LSmitll_NDROT-IN X42-LSmitll_SPLITT-OUT-X85-LSmitll_NDROT-IN X429-LSmitll_SPLITT-OUT-X85-LSmitll_NDROT-IN X85-LSmitll_NDROT-OUT-X87-LSmitll_SPLITT-INt LSmitll_NDROT

t992 X86-LSmitll_AND2T-OUT-X85-LSmitll_NDROT-INt 0 X86-LSmitll_AND2T-OUT-X85-LSmitll_NDROT-IN 0 z0=5 td=5.4ps
X86 X42-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-IN X83-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-IN X428-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-IN X86-LSmitll_AND2T-OUT-X85-LSmitll_NDROT-INt LSmitll_AND2T

t993 X87-LSmitll_SPLITT-OUT-X119-LSmitll_DFFT-INt 0 X87-LSmitll_SPLITT-OUT-X119-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t994 X87-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-INt 0 X87-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-IN 0 z0=5 td=1.1ps
X87 X85-LSmitll_NDROT-OUT-X87-LSmitll_SPLITT-IN X87-LSmitll_SPLITT-OUT-X119-LSmitll_DFFT-INt X87-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-INt LSmitll_SPLITT

t995 X88-LSmitll_NDROT-OUT-X90-LSmitll_SPLITT-INt 0 X88-LSmitll_NDROT-OUT-X90-LSmitll_SPLITT-IN 0 z0=5 td=12.4ps
X88 X89-LSmitll_AND2T-OUT-X88-LSmitll_NDROT-IN X43-LSmitll_SPLITT-OUT-X88-LSmitll_NDROT-IN X436-LSmitll_SPLITT-OUT-X88-LSmitll_NDROT-IN X88-LSmitll_NDROT-OUT-X90-LSmitll_SPLITT-INt LSmitll_NDROT

t996 X89-LSmitll_AND2T-OUT-X88-LSmitll_NDROT-INt 0 X89-LSmitll_AND2T-OUT-X88-LSmitll_NDROT-IN 0 z0=5 td=3.5ps
X89 X43-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-IN X84-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-IN X434-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-IN X89-LSmitll_AND2T-OUT-X88-LSmitll_NDROT-INt LSmitll_AND2T

t997 X90-LSmitll_SPLITT-OUT-X121-LSmitll_DFFT-INt 0 X90-LSmitll_SPLITT-OUT-X121-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t998 X90-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt 0 X90-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN 0 z0=5 td=5.9ps
X90 X88-LSmitll_NDROT-OUT-X90-LSmitll_SPLITT-IN X90-LSmitll_SPLITT-OUT-X121-LSmitll_DFFT-INt X90-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt LSmitll_SPLITT

t999 X91-LSmitll_NDROT-OUT-X93-LSmitll_SPLITT-INt 0 X91-LSmitll_NDROT-OUT-X93-LSmitll_SPLITT-IN 0 z0=5 td=10.5ps
X91 X92-LSmitll_AND2T-OUT-X91-LSmitll_NDROT-IN X45-LSmitll_SPLITT-OUT-X91-LSmitll_NDROT-IN X424-LSmitll_SPLITT-OUT-X91-LSmitll_NDROT-IN X91-LSmitll_NDROT-OUT-X93-LSmitll_SPLITT-INt LSmitll_NDROT

t1000 X92-LSmitll_AND2T-OUT-X91-LSmitll_NDROT-INt 0 X92-LSmitll_AND2T-OUT-X91-LSmitll_NDROT-IN 0 z0=5 td=3.4ps
X92 X45-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-IN X81-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-IN X429-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-IN X92-LSmitll_AND2T-OUT-X91-LSmitll_NDROT-INt LSmitll_AND2T

t1001 X93-LSmitll_SPLITT-OUT-X123-LSmitll_DFFT-INt 0 X93-LSmitll_SPLITT-OUT-X123-LSmitll_DFFT-IN 0 z0=5 td=5.7ps
t1002 X93-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt 0 X93-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X93 X91-LSmitll_NDROT-OUT-X93-LSmitll_SPLITT-IN X93-LSmitll_SPLITT-OUT-X123-LSmitll_DFFT-INt X93-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt LSmitll_SPLITT

t1003 X94-LSmitll_NDROT-OUT-X96-LSmitll_SPLITT-INt 0 X94-LSmitll_NDROT-OUT-X96-LSmitll_SPLITT-IN 0 z0=5 td=11.6ps
X94 X95-LSmitll_AND2T-OUT-X94-LSmitll_NDROT-IN X46-LSmitll_SPLITT-OUT-X94-LSmitll_NDROT-IN X527-LSmitll_SPLITT-OUT-X94-LSmitll_NDROT-IN X94-LSmitll_NDROT-OUT-X96-LSmitll_SPLITT-INt LSmitll_NDROT

t1004 X95-LSmitll_AND2T-OUT-X94-LSmitll_NDROT-INt 0 X95-LSmitll_AND2T-OUT-X94-LSmitll_NDROT-IN 0 z0=5 td=3.0ps
X95 X46-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-IN X82-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-IN X454-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-IN X95-LSmitll_AND2T-OUT-X94-LSmitll_NDROT-INt LSmitll_AND2T

t1005 X96-LSmitll_SPLITT-OUT-X125-LSmitll_DFFT-INt 0 X96-LSmitll_SPLITT-OUT-X125-LSmitll_DFFT-IN 0 z0=5 td=4.4ps
t1006 X96-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt 0 X96-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X96 X94-LSmitll_NDROT-OUT-X96-LSmitll_SPLITT-IN X96-LSmitll_SPLITT-OUT-X125-LSmitll_DFFT-INt X96-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt LSmitll_SPLITT

t1007 X97-LSmitll_NDROT-OUT-X99-LSmitll_SPLITT-INt 0 X97-LSmitll_NDROT-OUT-X99-LSmitll_SPLITT-IN 0 z0=5 td=7.7ps
X97 X98-LSmitll_AND2T-OUT-X97-LSmitll_NDROT-IN X48-LSmitll_SPLITT-OUT-X97-LSmitll_NDROT-IN X319-LSmitll_SPLITT-OUT-X97-LSmitll_NDROT-IN X97-LSmitll_NDROT-OUT-X99-LSmitll_SPLITT-INt LSmitll_NDROT

t1008 X98-LSmitll_AND2T-OUT-X97-LSmitll_NDROT-INt 0 X98-LSmitll_AND2T-OUT-X97-LSmitll_NDROT-IN 0 z0=5 td=1.4ps
X98 X48-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-IN X83-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-IN X528-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-IN X98-LSmitll_AND2T-OUT-X97-LSmitll_NDROT-INt LSmitll_AND2T

t1009 X99-LSmitll_SPLITT-OUT-X127-LSmitll_DFFT-INt 0 X99-LSmitll_SPLITT-OUT-X127-LSmitll_DFFT-IN 0 z0=5 td=4.1ps
t1010 X99-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt 0 X99-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN 0 z0=5 td=1.1ps
X99 X97-LSmitll_NDROT-OUT-X99-LSmitll_SPLITT-IN X99-LSmitll_SPLITT-OUT-X127-LSmitll_DFFT-INt X99-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt LSmitll_SPLITT

t1011 X100-LSmitll_NDROT-OUT-X102-LSmitll_SPLITT-INt 0 X100-LSmitll_NDROT-OUT-X102-LSmitll_SPLITT-IN 0 z0=5 td=12.6ps
X100 X101-LSmitll_AND2T-OUT-X100-LSmitll_NDROT-IN X49-LSmitll_SPLITT-OUT-X100-LSmitll_NDROT-IN X324-LSmitll_SPLITT-OUT-X100-LSmitll_NDROT-IN X100-LSmitll_NDROT-OUT-X102-LSmitll_SPLITT-INt LSmitll_NDROT

t1012 X101-LSmitll_AND2T-OUT-X100-LSmitll_NDROT-INt 0 X101-LSmitll_AND2T-OUT-X100-LSmitll_NDROT-IN 0 z0=5 td=2.6ps
X101 X49-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN X84-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN X324-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN X101-LSmitll_AND2T-OUT-X100-LSmitll_NDROT-INt LSmitll_AND2T

t1013 X102-LSmitll_SPLITT-OUT-X129-LSmitll_DFFT-INt 0 X102-LSmitll_SPLITT-OUT-X129-LSmitll_DFFT-IN 0 z0=5 td=2.9ps
t1014 X102-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-INt 0 X102-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X102 X100-LSmitll_NDROT-OUT-X102-LSmitll_SPLITT-IN X102-LSmitll_SPLITT-OUT-X129-LSmitll_DFFT-INt X102-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-INt LSmitll_SPLITT

t1015 X103-LSmitll_NDROT-OUT-X105-LSmitll_SPLITT-INt 0 X103-LSmitll_NDROT-OUT-X105-LSmitll_SPLITT-IN 0 z0=5 td=7.7ps
X103 X104-LSmitll_AND2T-OUT-X103-LSmitll_NDROT-IN X51-LSmitll_SPLITT-OUT-X103-LSmitll_NDROT-IN X319-LSmitll_SPLITT-OUT-X103-LSmitll_NDROT-IN X103-LSmitll_NDROT-OUT-X105-LSmitll_SPLITT-INt LSmitll_NDROT

t1016 X104-LSmitll_AND2T-OUT-X103-LSmitll_NDROT-INt 0 X104-LSmitll_AND2T-OUT-X103-LSmitll_NDROT-IN 0 z0=5 td=1.4ps
X104 X51-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN X81-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN X529-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN X104-LSmitll_AND2T-OUT-X103-LSmitll_NDROT-INt LSmitll_AND2T

t1017 X105-LSmitll_SPLITT-OUT-X131-LSmitll_DFFT-INt 0 X105-LSmitll_SPLITT-OUT-X131-LSmitll_DFFT-IN 0 z0=5 td=3.4ps
t1018 X105-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt 0 X105-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN 0 z0=5 td=6.0ps
X105 X103-LSmitll_NDROT-OUT-X105-LSmitll_SPLITT-IN X105-LSmitll_SPLITT-OUT-X131-LSmitll_DFFT-INt X105-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt LSmitll_SPLITT

t1019 X106-LSmitll_NDROT-OUT-X108-LSmitll_SPLITT-INt 0 X106-LSmitll_NDROT-OUT-X108-LSmitll_SPLITT-IN 0 z0=5 td=14.6ps
X106 X107-LSmitll_AND2T-OUT-X106-LSmitll_NDROT-IN X52-LSmitll_SPLITT-OUT-X106-LSmitll_NDROT-IN X530-LSmitll_SPLITT-OUT-X106-LSmitll_NDROT-IN X106-LSmitll_NDROT-OUT-X108-LSmitll_SPLITT-INt LSmitll_NDROT

t1020 X107-LSmitll_AND2T-OUT-X106-LSmitll_NDROT-INt 0 X107-LSmitll_AND2T-OUT-X106-LSmitll_NDROT-IN 0 z0=5 td=3.4ps
X107 X52-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN X82-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN X339-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN X107-LSmitll_AND2T-OUT-X106-LSmitll_NDROT-INt LSmitll_AND2T

t1021 X108-LSmitll_SPLITT-OUT-X133-LSmitll_DFFT-INt 0 X108-LSmitll_SPLITT-OUT-X133-LSmitll_DFFT-IN 0 z0=5 td=2.7ps
t1022 X108-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt 0 X108-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN 0 z0=5 td=1.1ps
X108 X106-LSmitll_NDROT-OUT-X108-LSmitll_SPLITT-IN X108-LSmitll_SPLITT-OUT-X133-LSmitll_DFFT-INt X108-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt LSmitll_SPLITT

t1023 X109-LSmitll_NDROT-OUT-X111-LSmitll_SPLITT-INt 0 X109-LSmitll_NDROT-OUT-X111-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X109 X110-LSmitll_AND2T-OUT-X109-LSmitll_NDROT-IN X55-LSmitll_SPLITT-OUT-X109-LSmitll_NDROT-IN X500-LSmitll_SPLITT-OUT-X109-LSmitll_NDROT-IN X109-LSmitll_NDROT-OUT-X111-LSmitll_SPLITT-INt LSmitll_NDROT

t1024 X110-LSmitll_AND2T-OUT-X109-LSmitll_NDROT-INt 0 X110-LSmitll_AND2T-OUT-X109-LSmitll_NDROT-IN 0 z0=5 td=3.0ps
X110 X55-LSmitll_SPLITT-OUT-X110-LSmitll_AND2T-IN X307-LSmitll_DFFT-OUT-X110-LSmitll_AND2T-IN X498-LSmitll_SPLITT-OUT-X110-LSmitll_AND2T-IN X110-LSmitll_AND2T-OUT-X109-LSmitll_NDROT-INt LSmitll_AND2T

t1025 X111-LSmitll_SPLITT-OUT-X135-LSmitll_DFFT-INt 0 X111-LSmitll_SPLITT-OUT-X135-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t1026 X111-LSmitll_SPLITT-OUT-X134-LSmitll_DFFT-INt 0 X111-LSmitll_SPLITT-OUT-X134-LSmitll_DFFT-IN 0 z0=5 td=8.7ps
X111 X109-LSmitll_NDROT-OUT-X111-LSmitll_SPLITT-IN X111-LSmitll_SPLITT-OUT-X135-LSmitll_DFFT-INt X111-LSmitll_SPLITT-OUT-X134-LSmitll_DFFT-INt LSmitll_SPLITT

t1027 X112-LSmitll_NDROT-OUT-X114-LSmitll_SPLITT-INt 0 X112-LSmitll_NDROT-OUT-X114-LSmitll_SPLITT-IN 0 z0=5 td=5.0ps
X112 X113-LSmitll_AND2T-OUT-X112-LSmitll_NDROT-IN X56-LSmitll_SPLITT-OUT-X112-LSmitll_NDROT-IN X475-LSmitll_SPLITT-OUT-X112-LSmitll_NDROT-IN X112-LSmitll_NDROT-OUT-X114-LSmitll_SPLITT-INt LSmitll_NDROT

t1028 X113-LSmitll_AND2T-OUT-X112-LSmitll_NDROT-INt 0 X113-LSmitll_AND2T-OUT-X112-LSmitll_NDROT-IN 0 z0=5 td=1.4ps
X113 X56-LSmitll_SPLITT-OUT-X113-LSmitll_AND2T-IN X308-LSmitll_DFFT-OUT-X113-LSmitll_AND2T-IN X531-LSmitll_SPLITT-OUT-X113-LSmitll_AND2T-IN X113-LSmitll_AND2T-OUT-X112-LSmitll_NDROT-INt LSmitll_AND2T

t1029 X114-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-INt 0 X114-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1030 X114-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-INt 0 X114-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-IN 0 z0=5 td=3.1ps
X114 X112-LSmitll_NDROT-OUT-X114-LSmitll_SPLITT-IN X114-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-INt X114-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-INt LSmitll_SPLITT

t1031 X115-LSmitll_NDROT-OUT-X117-LSmitll_SPLITT-INt 0 X115-LSmitll_NDROT-OUT-X117-LSmitll_SPLITT-IN 0 z0=5 td=7.4ps
X115 X116-LSmitll_AND2T-OUT-X115-LSmitll_NDROT-IN X53-LSmitll_SPLITT-OUT-X115-LSmitll_NDROT-IN X418-LSmitll_SPLITT-OUT-X115-LSmitll_NDROT-IN X115-LSmitll_NDROT-OUT-X117-LSmitll_SPLITT-INt LSmitll_NDROT

t1032 X116-LSmitll_AND2T-OUT-X115-LSmitll_NDROT-INt 0 X116-LSmitll_AND2T-OUT-X115-LSmitll_NDROT-IN 0 z0=5 td=1.4ps
X116 X53-LSmitll_SPLITT-OUT-X116-LSmitll_AND2T-IN X309-LSmitll_DFFT-OUT-X116-LSmitll_AND2T-IN X418-LSmitll_SPLITT-OUT-X116-LSmitll_AND2T-IN X116-LSmitll_AND2T-OUT-X115-LSmitll_NDROT-INt LSmitll_AND2T

t1033 X117-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-INt 0 X117-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-IN 0 z0=5 td=4.7ps
t1034 X117-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-INt 0 X117-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-IN 0 z0=5 td=3.2ps
X117 X115-LSmitll_NDROT-OUT-X117-LSmitll_SPLITT-IN X117-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-INt X117-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-INt LSmitll_SPLITT

t1035 X118-LSmitll_AND2T-OUT-X140-LSmitll_DFFT-INt 0 X118-LSmitll_AND2T-OUT-X140-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
X118 X69-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-IN X87-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-IN X482-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-IN X118-LSmitll_AND2T-OUT-X140-LSmitll_DFFT-INt LSmitll_AND2T


X119 X87-LSmitll_SPLITT-OUT-X119-LSmitll_DFFT-IN X487-LSmitll_SPLITT-OUT-X119-LSmitll_DFFT-IN reg1_out0_padt LSmitll_DFFT

t1037 X120-LSmitll_AND2T-OUT-X142-LSmitll_DFFT-INt 0 X120-LSmitll_AND2T-OUT-X142-LSmitll_DFFT-IN 0 z0=5 td=13.0ps
X120 X69-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN X90-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN X532-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN X120-LSmitll_AND2T-OUT-X142-LSmitll_DFFT-INt LSmitll_AND2T


X121 X90-LSmitll_SPLITT-OUT-X121-LSmitll_DFFT-IN X533-LSmitll_SPLITT-OUT-X121-LSmitll_DFFT-IN reg1_out1_padt LSmitll_DFFT

t1039 X122-LSmitll_AND2T-OUT-X144-LSmitll_DFFT-INt 0 X122-LSmitll_AND2T-OUT-X144-LSmitll_DFFT-IN 0 z0=5 td=2.4ps
X122 X70-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN X93-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN X504-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN X122-LSmitll_AND2T-OUT-X144-LSmitll_DFFT-INt LSmitll_AND2T


X123 X93-LSmitll_SPLITT-OUT-X123-LSmitll_DFFT-IN X408-LSmitll_SPLITT-OUT-X123-LSmitll_DFFT-IN reg1_out2_padt LSmitll_DFFT

t1041 X124-LSmitll_AND2T-OUT-X146-LSmitll_DFFT-INt 0 X124-LSmitll_AND2T-OUT-X146-LSmitll_DFFT-IN 0 z0=5 td=2.4ps
X124 X70-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN X96-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN X510-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN X124-LSmitll_AND2T-OUT-X146-LSmitll_DFFT-INt LSmitll_AND2T


X125 X96-LSmitll_SPLITT-OUT-X125-LSmitll_DFFT-IN X403-LSmitll_SPLITT-OUT-X125-LSmitll_DFFT-IN reg1_out3_padt LSmitll_DFFT

t1043 X126-LSmitll_AND2T-OUT-X141-LSmitll_XORT-INt 0 X126-LSmitll_AND2T-OUT-X141-LSmitll_XORT-IN 0 z0=5 td=4.0ps
X126 X71-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN X99-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN X381-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN X126-LSmitll_AND2T-OUT-X141-LSmitll_XORT-INt LSmitll_AND2T


X127 X99-LSmitll_SPLITT-OUT-X127-LSmitll_DFFT-IN X383-LSmitll_SPLITT-OUT-X127-LSmitll_DFFT-IN reg2_out0_padt LSmitll_DFFT

t1045 X128-LSmitll_AND2T-OUT-X143-LSmitll_XORT-INt 0 X128-LSmitll_AND2T-OUT-X143-LSmitll_XORT-IN 0 z0=5 td=2.8ps
X128 X71-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-IN X102-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-IN X376-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-IN X128-LSmitll_AND2T-OUT-X143-LSmitll_XORT-INt LSmitll_AND2T


X129 X102-LSmitll_SPLITT-OUT-X129-LSmitll_DFFT-IN X378-LSmitll_SPLITT-OUT-X129-LSmitll_DFFT-IN reg2_out1_padt LSmitll_DFFT

t1047 X130-LSmitll_AND2T-OUT-X145-LSmitll_XORT-INt 0 X130-LSmitll_AND2T-OUT-X145-LSmitll_XORT-IN 0 z0=5 td=4.0ps
X130 X72-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN X105-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN X534-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN X130-LSmitll_AND2T-OUT-X145-LSmitll_XORT-INt LSmitll_AND2T


X131 X105-LSmitll_SPLITT-OUT-X131-LSmitll_DFFT-IN X378-LSmitll_SPLITT-OUT-X131-LSmitll_DFFT-IN reg2_out2_padt LSmitll_DFFT

t1049 X132-LSmitll_AND2T-OUT-X147-LSmitll_XORT-INt 0 X132-LSmitll_AND2T-OUT-X147-LSmitll_XORT-IN 0 z0=5 td=4.4ps
X132 X72-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN X108-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN X480-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN X132-LSmitll_AND2T-OUT-X147-LSmitll_XORT-INt LSmitll_AND2T


X133 X108-LSmitll_SPLITT-OUT-X133-LSmitll_DFFT-IN X535-LSmitll_SPLITT-OUT-X133-LSmitll_DFFT-IN reg2_out3_padt LSmitll_DFFT


X134 X111-LSmitll_SPLITT-OUT-X134-LSmitll_DFFT-IN X536-LSmitll_SPLITT-OUT-X134-LSmitll_DFFT-IN regFlags_out0t LSmitll_DFFT


X135 X111-LSmitll_SPLITT-OUT-X135-LSmitll_DFFT-IN X537-LSmitll_SPLITT-OUT-X135-LSmitll_DFFT-IN regFlags_out0_padt LSmitll_DFFT


X136 X114-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-IN X538-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-IN regFlags_out1_padt LSmitll_DFFT


X137 X114-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-IN X507-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-IN regFlags_out1t LSmitll_DFFT


X138 X117-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-IN X539-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-IN regFlags_out2t LSmitll_DFFT


X139 X117-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-IN X449-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-IN regFlags_out2_padt LSmitll_DFFT

t1057 X140-LSmitll_DFFT-OUT-X149-LSmitll_SPLITT-INt 0 X140-LSmitll_DFFT-OUT-X149-LSmitll_SPLITT-IN 0 z0=5 td=8.1ps
X140 X118-LSmitll_AND2T-OUT-X140-LSmitll_DFFT-IN X482-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-IN X140-LSmitll_DFFT-OUT-X149-LSmitll_SPLITT-INt LSmitll_DFFT

t1058 X141-LSmitll_XORT-OUT-X148-LSmitll_SPLITT-INt 0 X141-LSmitll_XORT-OUT-X148-LSmitll_SPLITT-IN 0 z0=5 td=4.5ps
X141 X126-LSmitll_AND2T-OUT-X141-LSmitll_XORT-IN X17-LSmitll_SPLITT-OUT-X141-LSmitll_XORT-IN X400-LSmitll_SPLITT-OUT-X141-LSmitll_XORT-IN X141-LSmitll_XORT-OUT-X148-LSmitll_SPLITT-INt LSmitll_XORT

t1059 X142-LSmitll_DFFT-OUT-X151-LSmitll_SPLITT-INt 0 X142-LSmitll_DFFT-OUT-X151-LSmitll_SPLITT-IN 0 z0=5 td=6.0ps
X142 X120-LSmitll_AND2T-OUT-X142-LSmitll_DFFT-IN X383-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-IN X142-LSmitll_DFFT-OUT-X151-LSmitll_SPLITT-INt LSmitll_DFFT

t1060 X143-LSmitll_XORT-OUT-X150-LSmitll_SPLITT-INt 0 X143-LSmitll_XORT-OUT-X150-LSmitll_SPLITT-IN 0 z0=5 td=4.5ps
X143 X17-LSmitll_SPLITT-OUT-X143-LSmitll_XORT-IN X128-LSmitll_AND2T-OUT-X143-LSmitll_XORT-IN X540-LSmitll_SPLITT-OUT-X143-LSmitll_XORT-IN X143-LSmitll_XORT-OUT-X150-LSmitll_SPLITT-INt LSmitll_XORT

t1061 X144-LSmitll_DFFT-OUT-X153-LSmitll_SPLITT-INt 0 X144-LSmitll_DFFT-OUT-X153-LSmitll_SPLITT-IN 0 z0=5 td=6.0ps
X144 X122-LSmitll_AND2T-OUT-X144-LSmitll_DFFT-IN X505-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-IN X144-LSmitll_DFFT-OUT-X153-LSmitll_SPLITT-INt LSmitll_DFFT

t1062 X145-LSmitll_XORT-OUT-X152-LSmitll_SPLITT-INt 0 X145-LSmitll_XORT-OUT-X152-LSmitll_SPLITT-IN 0 z0=5 td=10.2ps
X145 X130-LSmitll_AND2T-OUT-X145-LSmitll_XORT-IN X18-LSmitll_SPLITT-OUT-X145-LSmitll_XORT-IN X479-LSmitll_SPLITT-OUT-X145-LSmitll_XORT-IN X145-LSmitll_XORT-OUT-X152-LSmitll_SPLITT-INt LSmitll_XORT

t1063 X146-LSmitll_DFFT-OUT-X155-LSmitll_SPLITT-INt 0 X146-LSmitll_DFFT-OUT-X155-LSmitll_SPLITT-IN 0 z0=5 td=14.2ps
X146 X124-LSmitll_AND2T-OUT-X146-LSmitll_DFFT-IN X512-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-IN X146-LSmitll_DFFT-OUT-X155-LSmitll_SPLITT-INt LSmitll_DFFT

t1064 X147-LSmitll_XORT-OUT-X154-LSmitll_SPLITT-INt 0 X147-LSmitll_XORT-OUT-X154-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X147 X18-LSmitll_SPLITT-OUT-X147-LSmitll_XORT-IN X132-LSmitll_AND2T-OUT-X147-LSmitll_XORT-IN X485-LSmitll_SPLITT-OUT-X147-LSmitll_XORT-IN X147-LSmitll_XORT-OUT-X154-LSmitll_SPLITT-INt LSmitll_XORT

t1065 X148-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-INt 0 X148-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-IN 0 z0=5 td=3.7ps
t1066 X148-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-INt 0 X148-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-IN 0 z0=5 td=1.9ps
X148 X141-LSmitll_XORT-OUT-X148-LSmitll_SPLITT-IN X148-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-INt X148-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-INt LSmitll_SPLITT

t1067 X149-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-INt 0 X149-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-IN 0 z0=5 td=1.9ps
t1068 X149-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-INt 0 X149-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-IN 0 z0=5 td=3.2ps
X149 X140-LSmitll_DFFT-OUT-X149-LSmitll_SPLITT-IN X149-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-INt X149-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-INt LSmitll_SPLITT

t1069 X150-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-INt 0 X150-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-IN 0 z0=5 td=4.9ps
t1070 X150-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-INt 0 X150-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-IN 0 z0=5 td=1.9ps
X150 X143-LSmitll_XORT-OUT-X150-LSmitll_SPLITT-IN X150-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-INt X150-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-INt LSmitll_SPLITT

t1071 X151-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-INt 0 X151-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-IN 0 z0=5 td=2.4ps
t1072 X151-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-INt 0 X151-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-IN 0 z0=5 td=1.1ps
X151 X142-LSmitll_DFFT-OUT-X151-LSmitll_SPLITT-IN X151-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-INt X151-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-INt LSmitll_SPLITT

t1073 X152-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-INt 0 X152-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-IN 0 z0=5 td=3.5ps
t1074 X152-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-INt 0 X152-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-IN 0 z0=5 td=3.9ps
X152 X145-LSmitll_XORT-OUT-X152-LSmitll_SPLITT-IN X152-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-INt X152-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-INt LSmitll_SPLITT

t1075 X153-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-INt 0 X153-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-IN 0 z0=5 td=2.5ps
t1076 X153-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-INt 0 X153-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-IN 0 z0=5 td=3.4ps
X153 X144-LSmitll_DFFT-OUT-X153-LSmitll_SPLITT-IN X153-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-INt X153-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-INt LSmitll_SPLITT

t1077 X154-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-INt 0 X154-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-IN 0 z0=5 td=3.7ps
t1078 X154-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-INt 0 X154-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-IN 0 z0=5 td=2.9ps
X154 X147-LSmitll_XORT-OUT-X154-LSmitll_SPLITT-IN X154-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-INt X154-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-INt LSmitll_SPLITT

t1079 X155-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-INt 0 X155-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-IN 0 z0=5 td=1.9ps
t1080 X155-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-INt 0 X155-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-IN 0 z0=5 td=2.8ps
X155 X146-LSmitll_DFFT-OUT-X155-LSmitll_SPLITT-IN X155-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-INt X155-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-INt LSmitll_SPLITT

t1081 X156-LSmitll_AND2T-OUT-X177-LSmitll_SPLITT-INt 0 X156-LSmitll_AND2T-OUT-X177-LSmitll_SPLITT-IN 0 z0=5 td=5.8ps
X156 X148-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-IN X149-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-IN X400-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-IN X156-LSmitll_AND2T-OUT-X177-LSmitll_SPLITT-INt LSmitll_AND2T

t1082 X157-LSmitll_XORT-OUT-X184-LSmitll_AND2T-INt 0 X157-LSmitll_XORT-OUT-X184-LSmitll_AND2T-IN 0 z0=5 td=11.7ps
X157 X148-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-IN X149-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-IN X401-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-IN X157-LSmitll_XORT-OUT-X184-LSmitll_AND2T-INt LSmitll_XORT

t1083 X158-LSmitll_AND2T-OUT-X178-LSmitll_SPLITT-INt 0 X158-LSmitll_AND2T-OUT-X178-LSmitll_SPLITT-IN 0 z0=5 td=10.1ps
X158 X150-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-IN X151-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-IN X381-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-IN X158-LSmitll_AND2T-OUT-X178-LSmitll_SPLITT-INt LSmitll_AND2T

t1084 X159-LSmitll_XORT-OUT-X187-LSmitll_AND2T-INt 0 X159-LSmitll_XORT-OUT-X187-LSmitll_AND2T-IN 0 z0=5 td=6.5ps
X159 X150-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-IN X151-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-IN X541-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-IN X159-LSmitll_XORT-OUT-X187-LSmitll_AND2T-INt LSmitll_XORT

t1085 X160-LSmitll_AND2T-OUT-X179-LSmitll_SPLITT-INt 0 X160-LSmitll_AND2T-OUT-X179-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X160 X152-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-IN X153-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-IN X500-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-IN X160-LSmitll_AND2T-OUT-X179-LSmitll_SPLITT-INt LSmitll_AND2T

t1086 X161-LSmitll_XORT-OUT-X190-LSmitll_AND2T-INt 0 X161-LSmitll_XORT-OUT-X190-LSmitll_AND2T-IN 0 z0=5 td=11.1ps
X161 X152-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-IN X153-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-IN X510-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-IN X161-LSmitll_XORT-OUT-X190-LSmitll_AND2T-INt LSmitll_XORT

t1087 X162-LSmitll_AND2T-OUT-X180-LSmitll_SPLITT-INt 0 X162-LSmitll_AND2T-OUT-X180-LSmitll_SPLITT-IN 0 z0=5 td=6.7ps
X162 X154-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-IN X155-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-IN X504-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-IN X162-LSmitll_AND2T-OUT-X180-LSmitll_SPLITT-INt LSmitll_AND2T

t1088 X163-LSmitll_XORT-OUT-X193-LSmitll_AND2T-INt 0 X163-LSmitll_XORT-OUT-X193-LSmitll_AND2T-IN 0 z0=5 td=10.5ps
X163 X154-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-IN X155-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-IN X505-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-IN X163-LSmitll_XORT-OUT-X193-LSmitll_AND2T-INt LSmitll_XORT

t1089 X164-LSmitll_DFFT-OUT-X168-LSmitll_SPLITT-INt 0 X164-LSmitll_DFFT-OUT-X168-LSmitll_SPLITT-IN 0 z0=5 td=8.1ps
X164 X20-LSmitll_DFFT-OUT-X164-LSmitll_DFFT-IN X323-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-IN X164-LSmitll_DFFT-OUT-X168-LSmitll_SPLITT-INt LSmitll_DFFT

t1090 X165-LSmitll_DFFT-OUT-X171-LSmitll_SPLITT-INt 0 X165-LSmitll_DFFT-OUT-X171-LSmitll_SPLITT-IN 0 z0=5 td=7.5ps
X165 X21-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-IN X512-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-IN X165-LSmitll_DFFT-OUT-X171-LSmitll_SPLITT-INt LSmitll_DFFT

t1091 X166-LSmitll_DFFT-OUT-X174-LSmitll_SPLITT-INt 0 X166-LSmitll_DFFT-OUT-X174-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
X166 X22-LSmitll_DFFT-OUT-X166-LSmitll_DFFT-IN X375-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-IN X166-LSmitll_DFFT-OUT-X174-LSmitll_SPLITT-INt LSmitll_DFFT

t1092 X167-LSmitll_DFFT-OUT-X181-LSmitll_DFFT-INt 0 X167-LSmitll_DFFT-OUT-X181-LSmitll_DFFT-IN 0 z0=5 td=5.2ps
X167 X19-LSmitll_DFFT-OUT-X167-LSmitll_DFFT-IN X363-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-IN X167-LSmitll_DFFT-OUT-X181-LSmitll_DFFT-INt LSmitll_DFFT

t1093 X168-LSmitll_SPLITT-OUT-X170-LSmitll_SPLITT-INt 0 X168-LSmitll_SPLITT-OUT-X170-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1094 X168-LSmitll_SPLITT-OUT-X169-LSmitll_SPLITT-INt 0 X168-LSmitll_SPLITT-OUT-X169-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X168 X164-LSmitll_DFFT-OUT-X168-LSmitll_SPLITT-IN X168-LSmitll_SPLITT-OUT-X170-LSmitll_SPLITT-INt X168-LSmitll_SPLITT-OUT-X169-LSmitll_SPLITT-INt LSmitll_SPLITT

t1095 X169-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-INt 0 X169-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1096 X169-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-INt 0 X169-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-IN 0 z0=5 td=4.1ps
X169 X168-LSmitll_SPLITT-OUT-X169-LSmitll_SPLITT-IN X169-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-INt X169-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-INt LSmitll_SPLITT

t1097 X170-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-INt 0 X170-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1098 X170-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-INt 0 X170-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-IN 0 z0=5 td=3.9ps
X170 X168-LSmitll_SPLITT-OUT-X170-LSmitll_SPLITT-IN X170-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-INt X170-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-INt LSmitll_SPLITT

t1099 X171-LSmitll_SPLITT-OUT-X173-LSmitll_SPLITT-INt 0 X171-LSmitll_SPLITT-OUT-X173-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
t1100 X171-LSmitll_SPLITT-OUT-X172-LSmitll_SPLITT-INt 0 X171-LSmitll_SPLITT-OUT-X172-LSmitll_SPLITT-IN 0 z0=5 td=4.9ps
X171 X165-LSmitll_DFFT-OUT-X171-LSmitll_SPLITT-IN X171-LSmitll_SPLITT-OUT-X173-LSmitll_SPLITT-INt X171-LSmitll_SPLITT-OUT-X172-LSmitll_SPLITT-INt LSmitll_SPLITT

t1101 X172-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-INt 0 X172-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-IN 0 z0=5 td=6.5ps
t1102 X172-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-INt 0 X172-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-IN 0 z0=5 td=1.1ps
X172 X171-LSmitll_SPLITT-OUT-X172-LSmitll_SPLITT-IN X172-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-INt X172-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-INt LSmitll_SPLITT

t1103 X173-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-INt 0 X173-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-IN 0 z0=5 td=4.9ps
t1104 X173-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-INt 0 X173-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-IN 0 z0=5 td=1.1ps
X173 X171-LSmitll_SPLITT-OUT-X173-LSmitll_SPLITT-IN X173-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-INt X173-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-INt LSmitll_SPLITT

t1105 X174-LSmitll_SPLITT-OUT-X176-LSmitll_SPLITT-INt 0 X174-LSmitll_SPLITT-OUT-X176-LSmitll_SPLITT-IN 0 z0=5 td=4.4ps
t1106 X174-LSmitll_SPLITT-OUT-X175-LSmitll_SPLITT-INt 0 X174-LSmitll_SPLITT-OUT-X175-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
X174 X166-LSmitll_DFFT-OUT-X174-LSmitll_SPLITT-IN X174-LSmitll_SPLITT-OUT-X176-LSmitll_SPLITT-INt X174-LSmitll_SPLITT-OUT-X175-LSmitll_SPLITT-INt LSmitll_SPLITT

t1107 X175-LSmitll_SPLITT-OUT-X187-LSmitll_AND2T-INt 0 X175-LSmitll_SPLITT-OUT-X187-LSmitll_AND2T-IN 0 z0=5 td=1.3ps
t1108 X175-LSmitll_SPLITT-OUT-X184-LSmitll_AND2T-INt 0 X175-LSmitll_SPLITT-OUT-X184-LSmitll_AND2T-IN 0 z0=5 td=5.3ps
X175 X174-LSmitll_SPLITT-OUT-X175-LSmitll_SPLITT-IN X175-LSmitll_SPLITT-OUT-X187-LSmitll_AND2T-INt X175-LSmitll_SPLITT-OUT-X184-LSmitll_AND2T-INt LSmitll_SPLITT

t1109 X176-LSmitll_SPLITT-OUT-X193-LSmitll_AND2T-INt 0 X176-LSmitll_SPLITT-OUT-X193-LSmitll_AND2T-IN 0 z0=5 td=3.5ps
t1110 X176-LSmitll_SPLITT-OUT-X190-LSmitll_AND2T-INt 0 X176-LSmitll_SPLITT-OUT-X190-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
X176 X174-LSmitll_SPLITT-OUT-X176-LSmitll_SPLITT-IN X176-LSmitll_SPLITT-OUT-X193-LSmitll_AND2T-INt X176-LSmitll_SPLITT-OUT-X190-LSmitll_AND2T-INt LSmitll_SPLITT

t1111 X177-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-INt 0 X177-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-IN 0 z0=5 td=3.2ps
t1112 X177-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-INt 0 X177-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-IN 0 z0=5 td=3.1ps
X177 X156-LSmitll_AND2T-OUT-X177-LSmitll_SPLITT-IN X177-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-INt X177-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-INt LSmitll_SPLITT

t1113 X178-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-INt 0 X178-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
t1114 X178-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-INt 0 X178-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-IN 0 z0=5 td=3.4ps
X178 X158-LSmitll_AND2T-OUT-X178-LSmitll_SPLITT-IN X178-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-INt X178-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-INt LSmitll_SPLITT

t1115 X179-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-INt 0 X179-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-IN 0 z0=5 td=3.6ps
t1116 X179-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-INt 0 X179-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-IN 0 z0=5 td=4.1ps
X179 X160-LSmitll_AND2T-OUT-X179-LSmitll_SPLITT-IN X179-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-INt X179-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-INt LSmitll_SPLITT

t1117 X180-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-INt 0 X180-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t1118 X180-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-INt 0 X180-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
X180 X162-LSmitll_AND2T-OUT-X180-LSmitll_SPLITT-IN X180-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-INt X180-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-INt LSmitll_SPLITT

t1119 X181-LSmitll_DFFT-OUT-X198-LSmitll_DFFT-INt 0 X181-LSmitll_DFFT-OUT-X198-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X181 X167-LSmitll_DFFT-OUT-X181-LSmitll_DFFT-IN X362-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-IN X181-LSmitll_DFFT-OUT-X198-LSmitll_DFFT-INt LSmitll_DFFT

t1120 X182-LSmitll_AND2T-OUT-X199-LSmitll_DFFT-INt 0 X182-LSmitll_AND2T-OUT-X199-LSmitll_DFFT-IN 0 z0=5 td=8.3ps
X182 X169-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-IN X177-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-IN X371-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-IN X182-LSmitll_AND2T-OUT-X199-LSmitll_DFFT-INt LSmitll_AND2T

t1121 X183-LSmitll_AND2T-OUT-X200-LSmitll_OR2T-INt 0 X183-LSmitll_AND2T-OUT-X200-LSmitll_OR2T-IN 0 z0=5 td=3.8ps
X183 X177-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-IN X172-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-IN X401-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-IN X183-LSmitll_AND2T-OUT-X200-LSmitll_OR2T-INt LSmitll_AND2T

t1122 X184-LSmitll_AND2T-OUT-X200-LSmitll_OR2T-INt 0 X184-LSmitll_AND2T-OUT-X200-LSmitll_OR2T-IN 0 z0=5 td=6.1ps
X184 X157-LSmitll_XORT-OUT-X184-LSmitll_AND2T-IN X175-LSmitll_SPLITT-OUT-X184-LSmitll_AND2T-IN X391-LSmitll_SPLITT-OUT-X184-LSmitll_AND2T-IN X184-LSmitll_AND2T-OUT-X200-LSmitll_OR2T-INt LSmitll_AND2T

t1123 X185-LSmitll_AND2T-OUT-X201-LSmitll_DFFT-INt 0 X185-LSmitll_AND2T-OUT-X201-LSmitll_DFFT-IN 0 z0=5 td=4.7ps
X185 X169-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-IN X178-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-IN X542-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-IN X185-LSmitll_AND2T-OUT-X201-LSmitll_DFFT-INt LSmitll_AND2T

t1124 X186-LSmitll_AND2T-OUT-X194-LSmitll_SPLITT-INt 0 X186-LSmitll_AND2T-OUT-X194-LSmitll_SPLITT-IN 0 z0=5 td=6.4ps
X186 X172-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-IN X178-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-IN X371-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-IN X186-LSmitll_AND2T-OUT-X194-LSmitll_SPLITT-INt LSmitll_AND2T

t1125 X187-LSmitll_AND2T-OUT-X195-LSmitll_SPLITT-INt 0 X187-LSmitll_AND2T-OUT-X195-LSmitll_SPLITT-IN 0 z0=5 td=4.9ps
X187 X159-LSmitll_XORT-OUT-X187-LSmitll_AND2T-IN X175-LSmitll_SPLITT-OUT-X187-LSmitll_AND2T-IN X376-LSmitll_SPLITT-OUT-X187-LSmitll_AND2T-IN X187-LSmitll_AND2T-OUT-X195-LSmitll_SPLITT-INt LSmitll_AND2T

t1126 X188-LSmitll_AND2T-OUT-X203-LSmitll_DFFT-INt 0 X188-LSmitll_AND2T-OUT-X203-LSmitll_DFFT-IN 0 z0=5 td=2.4ps
X188 X170-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-IN X179-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-IN X470-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-IN X188-LSmitll_AND2T-OUT-X203-LSmitll_DFFT-INt LSmitll_AND2T

t1127 X189-LSmitll_AND2T-OUT-X196-LSmitll_SPLITT-INt 0 X189-LSmitll_AND2T-OUT-X196-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
X189 X179-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-IN X173-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-IN X495-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-IN X189-LSmitll_AND2T-OUT-X196-LSmitll_SPLITT-INt LSmitll_AND2T

t1128 X190-LSmitll_AND2T-OUT-X197-LSmitll_SPLITT-INt 0 X190-LSmitll_AND2T-OUT-X197-LSmitll_SPLITT-IN 0 z0=5 td=4.5ps
X190 X161-LSmitll_XORT-OUT-X190-LSmitll_AND2T-IN X176-LSmitll_SPLITT-OUT-X190-LSmitll_AND2T-IN X543-LSmitll_SPLITT-OUT-X190-LSmitll_AND2T-IN X190-LSmitll_AND2T-OUT-X197-LSmitll_SPLITT-INt LSmitll_AND2T

t1129 X191-LSmitll_AND2T-OUT-X205-LSmitll_DFFT-INt 0 X191-LSmitll_AND2T-OUT-X205-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X191 X170-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-IN X180-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-IN X396-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-IN X191-LSmitll_AND2T-OUT-X205-LSmitll_DFFT-INt LSmitll_AND2T

t1130 X192-LSmitll_AND2T-OUT-X206-LSmitll_OR2T-INt 0 X192-LSmitll_AND2T-OUT-X206-LSmitll_OR2T-IN 0 z0=5 td=4.3ps
X192 X173-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-IN X180-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-IN X485-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-IN X192-LSmitll_AND2T-OUT-X206-LSmitll_OR2T-INt LSmitll_AND2T

t1131 X193-LSmitll_AND2T-OUT-X206-LSmitll_OR2T-INt 0 X193-LSmitll_AND2T-OUT-X206-LSmitll_OR2T-IN 0 z0=5 td=1.4ps
X193 X163-LSmitll_XORT-OUT-X193-LSmitll_AND2T-IN X176-LSmitll_SPLITT-OUT-X193-LSmitll_AND2T-IN X479-LSmitll_SPLITT-OUT-X193-LSmitll_AND2T-IN X193-LSmitll_AND2T-OUT-X206-LSmitll_OR2T-INt LSmitll_AND2T

t1132 X194-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-INt 0 X194-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-IN 0 z0=5 td=1.3ps
t1133 X194-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-INt 0 X194-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-IN 0 z0=5 td=2.8ps
X194 X186-LSmitll_AND2T-OUT-X194-LSmitll_SPLITT-IN X194-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-INt X194-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-INt LSmitll_SPLITT

t1134 X195-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-INt 0 X195-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-IN 0 z0=5 td=3.9ps
t1135 X195-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-INt 0 X195-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-IN 0 z0=5 td=2.6ps
X195 X187-LSmitll_AND2T-OUT-X195-LSmitll_SPLITT-IN X195-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-INt X195-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-INt LSmitll_SPLITT

t1136 X196-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-INt 0 X196-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-IN 0 z0=5 td=3.6ps
t1137 X196-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-INt 0 X196-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-IN 0 z0=5 td=1.1ps
X196 X189-LSmitll_AND2T-OUT-X196-LSmitll_SPLITT-IN X196-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-INt X196-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-INt LSmitll_SPLITT

t1138 X197-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-INt 0 X197-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-IN 0 z0=5 td=1.9ps
t1139 X197-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-INt 0 X197-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-IN 0 z0=5 td=2.6ps
X197 X190-LSmitll_AND2T-OUT-X197-LSmitll_SPLITT-IN X197-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-INt X197-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-INt LSmitll_SPLITT

t1140 X198-LSmitll_DFFT-OUT-X224-LSmitll_SPLITT-INt 0 X198-LSmitll_DFFT-OUT-X224-LSmitll_SPLITT-IN 0 z0=5 td=11.6ps
X198 X181-LSmitll_DFFT-OUT-X198-LSmitll_DFFT-IN X326-LSmitll_SPLITT-OUT-X198-LSmitll_DFFT-IN X198-LSmitll_DFFT-OUT-X224-LSmitll_SPLITT-INt LSmitll_DFFT

t1141 X199-LSmitll_DFFT-OUT-X209-LSmitll_SPLITT-INt 0 X199-LSmitll_DFFT-OUT-X209-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X199 X182-LSmitll_AND2T-OUT-X199-LSmitll_DFFT-IN X363-LSmitll_SPLITT-OUT-X199-LSmitll_DFFT-IN X199-LSmitll_DFFT-OUT-X209-LSmitll_SPLITT-INt LSmitll_DFFT

t1142 X200-LSmitll_OR2T-OUT-X210-LSmitll_SPLITT-INt 0 X200-LSmitll_OR2T-OUT-X210-LSmitll_SPLITT-IN 0 z0=5 td=6.5ps
X200 X183-LSmitll_AND2T-OUT-X200-LSmitll_OR2T-IN X184-LSmitll_AND2T-OUT-X200-LSmitll_OR2T-IN X406-LSmitll_SPLITT-OUT-X200-LSmitll_OR2T-IN X200-LSmitll_OR2T-OUT-X210-LSmitll_SPLITT-INt LSmitll_OR2T

t1143 X201-LSmitll_DFFT-OUT-X213-LSmitll_SPLITT-INt 0 X201-LSmitll_DFFT-OUT-X213-LSmitll_SPLITT-IN 0 z0=5 td=9.7ps
X201 X185-LSmitll_AND2T-OUT-X201-LSmitll_DFFT-IN X365-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-IN X201-LSmitll_DFFT-OUT-X213-LSmitll_SPLITT-INt LSmitll_DFFT

t1144 X202-LSmitll_OR2T-OUT-X214-LSmitll_SPLITT-INt 0 X202-LSmitll_OR2T-OUT-X214-LSmitll_SPLITT-IN 0 z0=5 td=4.7ps
X202 X194-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-IN X195-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-IN X544-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-IN X202-LSmitll_OR2T-OUT-X214-LSmitll_SPLITT-INt LSmitll_OR2T

t1145 X203-LSmitll_DFFT-OUT-X217-LSmitll_SPLITT-INt 0 X203-LSmitll_DFFT-OUT-X217-LSmitll_SPLITT-IN 0 z0=5 td=6.2ps
X203 X188-LSmitll_AND2T-OUT-X203-LSmitll_DFFT-IN X470-LSmitll_SPLITT-OUT-X203-LSmitll_DFFT-IN X203-LSmitll_DFFT-OUT-X217-LSmitll_SPLITT-INt LSmitll_DFFT

t1146 X204-LSmitll_OR2T-OUT-X218-LSmitll_SPLITT-INt 0 X204-LSmitll_OR2T-OUT-X218-LSmitll_SPLITT-IN 0 z0=5 td=5.0ps
X204 X196-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-IN X197-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-IN X475-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-IN X204-LSmitll_OR2T-OUT-X218-LSmitll_SPLITT-INt LSmitll_OR2T

t1147 X205-LSmitll_DFFT-OUT-X236-LSmitll_DFFT-INt 0 X205-LSmitll_DFFT-OUT-X236-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X205 X191-LSmitll_AND2T-OUT-X205-LSmitll_DFFT-IN X396-LSmitll_SPLITT-OUT-X205-LSmitll_DFFT-IN X205-LSmitll_DFFT-OUT-X236-LSmitll_DFFT-INt LSmitll_DFFT

t1148 X206-LSmitll_OR2T-OUT-X221-LSmitll_SPLITT-INt 0 X206-LSmitll_OR2T-OUT-X221-LSmitll_SPLITT-IN 0 z0=5 td=8.8ps
X206 X192-LSmitll_AND2T-OUT-X206-LSmitll_OR2T-IN X193-LSmitll_AND2T-OUT-X206-LSmitll_OR2T-IN X545-LSmitll_SPLITT-OUT-X206-LSmitll_OR2T-IN X206-LSmitll_OR2T-OUT-X221-LSmitll_SPLITT-INt LSmitll_OR2T

t1149 X207-LSmitll_OR2T-OUT-X215-LSmitll_SPLITT-INt 0 X207-LSmitll_OR2T-OUT-X215-LSmitll_SPLITT-IN 0 z0=5 td=7.0ps
X207 X194-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-IN X195-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-IN X391-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-IN X207-LSmitll_OR2T-OUT-X215-LSmitll_SPLITT-INt LSmitll_OR2T

t1150 X208-LSmitll_OR2T-OUT-X219-LSmitll_SPLITT-INt 0 X208-LSmitll_OR2T-OUT-X219-LSmitll_SPLITT-IN 0 z0=5 td=14.3ps
X208 X196-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-IN X197-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-IN X480-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-IN X208-LSmitll_OR2T-OUT-X219-LSmitll_SPLITT-INt LSmitll_OR2T

t1151 X209-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-INt 0 X209-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1152 X209-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-INt 0 X209-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-IN 0 z0=5 td=4.7ps
X209 X199-LSmitll_DFFT-OUT-X209-LSmitll_SPLITT-IN X209-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-INt X209-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-INt LSmitll_SPLITT

t1153 X210-LSmitll_SPLITT-OUT-X212-LSmitll_SPLITT-INt 0 X210-LSmitll_SPLITT-OUT-X212-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1154 X210-LSmitll_SPLITT-OUT-X211-LSmitll_SPLITT-INt 0 X210-LSmitll_SPLITT-OUT-X211-LSmitll_SPLITT-IN 0 z0=5 td=8.4ps
X210 X200-LSmitll_OR2T-OUT-X210-LSmitll_SPLITT-IN X210-LSmitll_SPLITT-OUT-X212-LSmitll_SPLITT-INt X210-LSmitll_SPLITT-OUT-X211-LSmitll_SPLITT-INt LSmitll_SPLITT

t1155 X211-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-INt 0 X211-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-IN 0 z0=5 td=7.1ps
t1156 X211-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-INt 0 X211-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-IN 0 z0=5 td=2.0ps
X211 X210-LSmitll_SPLITT-OUT-X211-LSmitll_SPLITT-IN X211-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-INt X211-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-INt LSmitll_SPLITT

t1157 X212-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt 0 X212-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN 0 z0=5 td=7.8ps
t1158 X212-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-INt 0 X212-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-IN 0 z0=5 td=13.5ps
X212 X210-LSmitll_SPLITT-OUT-X212-LSmitll_SPLITT-IN X212-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt X212-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-INt LSmitll_SPLITT

t1159 X213-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt 0 X213-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN 0 z0=5 td=3.4ps
t1160 X213-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-INt 0 X213-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
X213 X201-LSmitll_DFFT-OUT-X213-LSmitll_SPLITT-IN X213-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt X213-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-INt LSmitll_SPLITT

t1161 X214-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-INt 0 X214-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-IN 0 z0=5 td=2.6ps
t1162 X214-LSmitll_SPLITT-OUT-X229-LSmitll_DFFT-INt 0 X214-LSmitll_SPLITT-OUT-X229-LSmitll_DFFT-IN 0 z0=5 td=6.1ps
X214 X202-LSmitll_OR2T-OUT-X214-LSmitll_SPLITT-IN X214-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-INt X214-LSmitll_SPLITT-OUT-X229-LSmitll_DFFT-INt LSmitll_SPLITT

t1163 X215-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt 0 X215-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN 0 z0=5 td=4.3ps
t1164 X215-LSmitll_SPLITT-OUT-X216-LSmitll_SPLITT-INt 0 X215-LSmitll_SPLITT-OUT-X216-LSmitll_SPLITT-IN 0 z0=5 td=8.2ps
X215 X207-LSmitll_OR2T-OUT-X215-LSmitll_SPLITT-IN X215-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt X215-LSmitll_SPLITT-OUT-X216-LSmitll_SPLITT-INt LSmitll_SPLITT

t1165 X216-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-INt 0 X216-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1166 X216-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-INt 0 X216-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-IN 0 z0=5 td=2.6ps
X216 X215-LSmitll_SPLITT-OUT-X216-LSmitll_SPLITT-IN X216-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-INt X216-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-INt LSmitll_SPLITT

t1167 X217-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt 0 X217-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN 0 z0=5 td=2.9ps
t1168 X217-LSmitll_SPLITT-OUT-X232-LSmitll_DFFT-INt 0 X217-LSmitll_SPLITT-OUT-X232-LSmitll_DFFT-IN 0 z0=5 td=4.4ps
X217 X203-LSmitll_DFFT-OUT-X217-LSmitll_SPLITT-IN X217-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt X217-LSmitll_SPLITT-OUT-X232-LSmitll_DFFT-INt LSmitll_SPLITT

t1169 X218-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt 0 X218-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t1170 X218-LSmitll_SPLITT-OUT-X233-LSmitll_DFFT-INt 0 X218-LSmitll_SPLITT-OUT-X233-LSmitll_DFFT-IN 0 z0=5 td=5.1ps
X218 X204-LSmitll_OR2T-OUT-X218-LSmitll_SPLITT-IN X218-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt X218-LSmitll_SPLITT-OUT-X233-LSmitll_DFFT-INt LSmitll_SPLITT

t1171 X219-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-INt 0 X219-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-IN 0 z0=5 td=1.3ps
t1172 X219-LSmitll_SPLITT-OUT-X220-LSmitll_SPLITT-INt 0 X219-LSmitll_SPLITT-OUT-X220-LSmitll_SPLITT-IN 0 z0=5 td=3.5ps
X219 X208-LSmitll_OR2T-OUT-X219-LSmitll_SPLITT-IN X219-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-INt X219-LSmitll_SPLITT-OUT-X220-LSmitll_SPLITT-INt LSmitll_SPLITT

t1173 X220-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-INt 0 X220-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-IN 0 z0=5 td=3.6ps
t1174 X220-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-INt 0 X220-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-IN 0 z0=5 td=3.3ps
X220 X219-LSmitll_SPLITT-OUT-X220-LSmitll_SPLITT-IN X220-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-INt X220-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-INt LSmitll_SPLITT

t1175 X221-LSmitll_SPLITT-OUT-X223-LSmitll_SPLITT-INt 0 X221-LSmitll_SPLITT-OUT-X223-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
t1176 X221-LSmitll_SPLITT-OUT-X222-LSmitll_SPLITT-INt 0 X221-LSmitll_SPLITT-OUT-X222-LSmitll_SPLITT-IN 0 z0=5 td=5.3ps
X221 X206-LSmitll_OR2T-OUT-X221-LSmitll_SPLITT-IN X221-LSmitll_SPLITT-OUT-X223-LSmitll_SPLITT-INt X221-LSmitll_SPLITT-OUT-X222-LSmitll_SPLITT-INt LSmitll_SPLITT

t1177 X222-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt 0 X222-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
t1178 X222-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-INt 0 X222-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-IN 0 z0=5 td=7.1ps
X222 X221-LSmitll_SPLITT-OUT-X222-LSmitll_SPLITT-IN X222-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt X222-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-INt LSmitll_SPLITT

t1179 X223-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-INt 0 X223-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-IN 0 z0=5 td=4.0ps
t1180 X223-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-INt 0 X223-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-IN 0 z0=5 td=6.3ps
X223 X221-LSmitll_SPLITT-OUT-X223-LSmitll_SPLITT-IN X223-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-INt X223-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-INt LSmitll_SPLITT

t1181 X224-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-INt 0 X224-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t1182 X224-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-INt 0 X224-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-IN 0 z0=5 td=6.7ps
X224 X198-LSmitll_DFFT-OUT-X224-LSmitll_SPLITT-IN X224-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-INt X224-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-INt LSmitll_SPLITT

t1183 X225-LSmitll_DFFT-OUT-X244-LSmitll_OR2T-INt 0 X225-LSmitll_DFFT-OUT-X244-LSmitll_OR2T-IN 0 z0=5 td=9.4ps
X225 X209-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-IN X546-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-IN X225-LSmitll_DFFT-OUT-X244-LSmitll_OR2T-INt LSmitll_DFFT

t1184 X226-LSmitll_DFFT-OUT-X243-LSmitll_DFFT-INt 0 X226-LSmitll_DFFT-OUT-X243-LSmitll_DFFT-IN 0 z0=5 td=10.9ps
X226 X211-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-IN X349-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-IN X226-LSmitll_DFFT-OUT-X243-LSmitll_DFFT-INt LSmitll_DFFT

t1185 X227-LSmitll_AND2T-OUT-X244-LSmitll_OR2T-INt 0 X227-LSmitll_AND2T-OUT-X244-LSmitll_OR2T-IN 0 z0=5 td=13.4ps
X227 X211-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-IN X224-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-IN X331-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-IN X227-LSmitll_AND2T-OUT-X244-LSmitll_OR2T-INt LSmitll_AND2T

t1186 X228-LSmitll_DFFT-OUT-X246-LSmitll_OR2T-INt 0 X228-LSmitll_DFFT-OUT-X246-LSmitll_OR2T-IN 0 z0=5 td=7.8ps
X228 X213-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-IN X388-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-IN X228-LSmitll_DFFT-OUT-X246-LSmitll_OR2T-INt LSmitll_DFFT

t1187 X229-LSmitll_DFFT-OUT-X245-LSmitll_DFFT-INt 0 X229-LSmitll_DFFT-OUT-X245-LSmitll_DFFT-IN 0 z0=5 td=14.8ps
X229 X214-LSmitll_SPLITT-OUT-X229-LSmitll_DFFT-IN X329-LSmitll_SPLITT-OUT-X229-LSmitll_DFFT-IN X229-LSmitll_DFFT-OUT-X245-LSmitll_DFFT-INt LSmitll_DFFT

t1188 X230-LSmitll_AND2T-OUT-X246-LSmitll_OR2T-INt 0 X230-LSmitll_AND2T-OUT-X246-LSmitll_OR2T-IN 0 z0=5 td=5.9ps
X230 X209-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-IN X214-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-IN X368-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-IN X230-LSmitll_AND2T-OUT-X246-LSmitll_OR2T-INt LSmitll_AND2T

t1189 X231-LSmitll_AND2T-OUT-X247-LSmitll_DFFT-INt 0 X231-LSmitll_AND2T-OUT-X247-LSmitll_DFFT-IN 0 z0=5 td=14.5ps
X231 X212-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-IN X216-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-IN X467-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-IN X231-LSmitll_AND2T-OUT-X247-LSmitll_DFFT-INt LSmitll_AND2T

t1190 X232-LSmitll_DFFT-OUT-X249-LSmitll_OR2T-INt 0 X232-LSmitll_DFFT-OUT-X249-LSmitll_OR2T-IN 0 z0=5 td=1.0ps
X232 X217-LSmitll_SPLITT-OUT-X232-LSmitll_DFFT-IN X493-LSmitll_SPLITT-OUT-X232-LSmitll_DFFT-IN X232-LSmitll_DFFT-OUT-X249-LSmitll_OR2T-INt LSmitll_DFFT

t1191 X233-LSmitll_DFFT-OUT-X248-LSmitll_DFFT-INt 0 X233-LSmitll_DFFT-OUT-X248-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X233 X218-LSmitll_SPLITT-OUT-X233-LSmitll_DFFT-IN X436-LSmitll_SPLITT-OUT-X233-LSmitll_DFFT-IN X233-LSmitll_DFFT-OUT-X248-LSmitll_DFFT-INt LSmitll_DFFT

t1192 X234-LSmitll_AND2T-OUT-X249-LSmitll_OR2T-INt 0 X234-LSmitll_AND2T-OUT-X249-LSmitll_OR2T-IN 0 z0=5 td=2.8ps
X234 X213-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN X218-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN X492-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN X234-LSmitll_AND2T-OUT-X249-LSmitll_OR2T-INt LSmitll_AND2T

t1193 X235-LSmitll_AND2T-OUT-X250-LSmitll_DFFT-INt 0 X235-LSmitll_AND2T-OUT-X250-LSmitll_DFFT-IN 0 z0=5 td=2.4ps
X235 X216-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-IN X220-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-IN X468-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-IN X235-LSmitll_AND2T-OUT-X250-LSmitll_DFFT-INt LSmitll_AND2T

t1194 X236-LSmitll_DFFT-OUT-X252-LSmitll_OR2T-INt 0 X236-LSmitll_DFFT-OUT-X252-LSmitll_OR2T-IN 0 z0=5 td=3.9ps
X236 X205-LSmitll_DFFT-OUT-X236-LSmitll_DFFT-IN X547-LSmitll_SPLITT-OUT-X236-LSmitll_DFFT-IN X236-LSmitll_DFFT-OUT-X252-LSmitll_OR2T-INt LSmitll_DFFT

t1195 X237-LSmitll_DFFT-OUT-X251-LSmitll_DFFT-INt 0 X237-LSmitll_DFFT-OUT-X251-LSmitll_DFFT-IN 0 z0=5 td=9.5ps
X237 X222-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-IN X498-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-IN X237-LSmitll_DFFT-OUT-X251-LSmitll_DFFT-INt LSmitll_DFFT

t1196 X238-LSmitll_AND2T-OUT-X252-LSmitll_OR2T-INt 0 X238-LSmitll_AND2T-OUT-X252-LSmitll_OR2T-IN 0 z0=5 td=1.4ps
X238 X217-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN X222-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN X394-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN X238-LSmitll_AND2T-OUT-X252-LSmitll_OR2T-INt LSmitll_AND2T

t1197 X239-LSmitll_AND2T-OUT-X253-LSmitll_DFFT-INt 0 X239-LSmitll_AND2T-OUT-X253-LSmitll_DFFT-IN 0 z0=5 td=2.4ps
X239 X220-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-IN X223-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-IN X388-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-IN X239-LSmitll_AND2T-OUT-X253-LSmitll_DFFT-INt LSmitll_AND2T

t1198 X240-LSmitll_AND2T-OUT-X254-LSmitll_AND2T-INt 0 X240-LSmitll_AND2T-OUT-X254-LSmitll_AND2T-IN 0 z0=5 td=2.6ps
X240 X212-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN X215-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN X365-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN X240-LSmitll_AND2T-OUT-X254-LSmitll_AND2T-INt LSmitll_AND2T

t1199 X241-LSmitll_AND2T-OUT-X254-LSmitll_AND2T-INt 0 X241-LSmitll_AND2T-OUT-X254-LSmitll_AND2T-IN 0 z0=5 td=10.2ps
X241 X219-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-IN X223-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-IN X369-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-IN X241-LSmitll_AND2T-OUT-X254-LSmitll_AND2T-INt LSmitll_AND2T

t1200 X242-LSmitll_DFFT-OUT-X255-LSmitll_DFFT-INt 0 X242-LSmitll_DFFT-OUT-X255-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X242 X224-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-IN X326-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-IN X242-LSmitll_DFFT-OUT-X255-LSmitll_DFFT-INt LSmitll_DFFT

t1201 X243-LSmitll_DFFT-OUT-X262-LSmitll_DFFT-INt 0 X243-LSmitll_DFFT-OUT-X262-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X243 X226-LSmitll_DFFT-OUT-X243-LSmitll_DFFT-IN X548-LSmitll_SPLITT-OUT-X243-LSmitll_DFFT-IN X243-LSmitll_DFFT-OUT-X262-LSmitll_DFFT-INt LSmitll_DFFT

t1202 X244-LSmitll_OR2T-OUT-X257-LSmitll_SPLITT-INt 0 X244-LSmitll_OR2T-OUT-X257-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X244 X225-LSmitll_DFFT-OUT-X244-LSmitll_OR2T-IN X227-LSmitll_AND2T-OUT-X244-LSmitll_OR2T-IN X549-LSmitll_SPLITT-OUT-X244-LSmitll_OR2T-IN X244-LSmitll_OR2T-OUT-X257-LSmitll_SPLITT-INt LSmitll_OR2T

t1203 X245-LSmitll_DFFT-OUT-X264-LSmitll_DFFT-INt 0 X245-LSmitll_DFFT-OUT-X264-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X245 X229-LSmitll_DFFT-OUT-X245-LSmitll_DFFT-IN X348-LSmitll_SPLITT-OUT-X245-LSmitll_DFFT-IN X245-LSmitll_DFFT-OUT-X264-LSmitll_DFFT-INt LSmitll_DFFT

t1204 X246-LSmitll_OR2T-OUT-X258-LSmitll_SPLITT-INt 0 X246-LSmitll_OR2T-OUT-X258-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X246 X228-LSmitll_DFFT-OUT-X246-LSmitll_OR2T-IN X230-LSmitll_AND2T-OUT-X246-LSmitll_OR2T-IN X331-LSmitll_SPLITT-OUT-X246-LSmitll_OR2T-IN X246-LSmitll_OR2T-OUT-X258-LSmitll_SPLITT-INt LSmitll_OR2T

t1205 X247-LSmitll_DFFT-OUT-X259-LSmitll_SPLITT-INt 0 X247-LSmitll_DFFT-OUT-X259-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X247 X231-LSmitll_AND2T-OUT-X247-LSmitll_DFFT-IN X351-LSmitll_SPLITT-OUT-X247-LSmitll_DFFT-IN X247-LSmitll_DFFT-OUT-X259-LSmitll_SPLITT-INt LSmitll_DFFT

t1206 X248-LSmitll_DFFT-OUT-X267-LSmitll_DFFT-INt 0 X248-LSmitll_DFFT-OUT-X267-LSmitll_DFFT-IN 0 z0=5 td=5.4ps
X248 X233-LSmitll_DFFT-OUT-X248-LSmitll_DFFT-IN X473-LSmitll_SPLITT-OUT-X248-LSmitll_DFFT-IN X248-LSmitll_DFFT-OUT-X267-LSmitll_DFFT-INt LSmitll_DFFT

t1207 X249-LSmitll_OR2T-OUT-X268-LSmitll_DFFT-INt 0 X249-LSmitll_OR2T-OUT-X268-LSmitll_DFFT-IN 0 z0=5 td=9.4ps
X249 X232-LSmitll_DFFT-OUT-X249-LSmitll_OR2T-IN X234-LSmitll_AND2T-OUT-X249-LSmitll_OR2T-IN X493-LSmitll_SPLITT-OUT-X249-LSmitll_OR2T-IN X249-LSmitll_OR2T-OUT-X268-LSmitll_DFFT-INt LSmitll_OR2T

t1208 X250-LSmitll_DFFT-OUT-X269-LSmitll_AND2T-INt 0 X250-LSmitll_DFFT-OUT-X269-LSmitll_AND2T-IN 0 z0=5 td=9.8ps
X250 X235-LSmitll_AND2T-OUT-X250-LSmitll_DFFT-IN X473-LSmitll_SPLITT-OUT-X250-LSmitll_DFFT-IN X250-LSmitll_DFFT-OUT-X269-LSmitll_AND2T-INt LSmitll_DFFT

t1209 X251-LSmitll_DFFT-OUT-X270-LSmitll_DFFT-INt 0 X251-LSmitll_DFFT-OUT-X270-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X251 X237-LSmitll_DFFT-OUT-X251-LSmitll_DFFT-IN X550-LSmitll_SPLITT-OUT-X251-LSmitll_DFFT-IN X251-LSmitll_DFFT-OUT-X270-LSmitll_DFFT-INt LSmitll_DFFT

t1210 X252-LSmitll_OR2T-OUT-X271-LSmitll_DFFT-INt 0 X252-LSmitll_OR2T-OUT-X271-LSmitll_DFFT-IN 0 z0=5 td=8.3ps
X252 X236-LSmitll_DFFT-OUT-X252-LSmitll_OR2T-IN X238-LSmitll_AND2T-OUT-X252-LSmitll_OR2T-IN X389-LSmitll_SPLITT-OUT-X252-LSmitll_OR2T-IN X252-LSmitll_OR2T-OUT-X271-LSmitll_DFFT-INt LSmitll_OR2T

t1211 X253-LSmitll_DFFT-OUT-X260-LSmitll_SPLITT-INt 0 X253-LSmitll_DFFT-OUT-X260-LSmitll_SPLITT-IN 0 z0=5 td=8.5ps
X253 X239-LSmitll_AND2T-OUT-X253-LSmitll_DFFT-IN X389-LSmitll_SPLITT-OUT-X253-LSmitll_DFFT-IN X253-LSmitll_DFFT-OUT-X260-LSmitll_SPLITT-INt LSmitll_DFFT

t1212 X254-LSmitll_AND2T-OUT-X274-LSmitll_DFFT-INt 0 X254-LSmitll_AND2T-OUT-X274-LSmitll_DFFT-IN 0 z0=5 td=5.1ps
X254 X240-LSmitll_AND2T-OUT-X254-LSmitll_AND2T-IN X241-LSmitll_AND2T-OUT-X254-LSmitll_AND2T-IN X368-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-IN X254-LSmitll_AND2T-OUT-X274-LSmitll_DFFT-INt LSmitll_AND2T

t1213 X255-LSmitll_DFFT-OUT-X256-LSmitll_SPLITT-INt 0 X255-LSmitll_DFFT-OUT-X256-LSmitll_SPLITT-IN 0 z0=5 td=13.1ps
X255 X242-LSmitll_DFFT-OUT-X255-LSmitll_DFFT-IN X329-LSmitll_SPLITT-OUT-X255-LSmitll_DFFT-IN X255-LSmitll_DFFT-OUT-X256-LSmitll_SPLITT-INt LSmitll_DFFT

t1214 X256-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt 0 X256-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1215 X256-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-INt 0 X256-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-IN 0 z0=5 td=7.4ps
X256 X255-LSmitll_DFFT-OUT-X256-LSmitll_SPLITT-IN X256-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt X256-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-INt LSmitll_SPLITT

t1216 X257-LSmitll_SPLITT-OUT-X269-LSmitll_AND2T-INt 0 X257-LSmitll_SPLITT-OUT-X269-LSmitll_AND2T-IN 0 z0=5 td=3.5ps
t1217 X257-LSmitll_SPLITT-OUT-X263-LSmitll_DFFT-INt 0 X257-LSmitll_SPLITT-OUT-X263-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
X257 X244-LSmitll_OR2T-OUT-X257-LSmitll_SPLITT-IN X257-LSmitll_SPLITT-OUT-X269-LSmitll_AND2T-INt X257-LSmitll_SPLITT-OUT-X263-LSmitll_DFFT-INt LSmitll_SPLITT

t1218 X258-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-INt 0 X258-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
t1219 X258-LSmitll_SPLITT-OUT-X265-LSmitll_DFFT-INt 0 X258-LSmitll_SPLITT-OUT-X265-LSmitll_DFFT-IN 0 z0=5 td=4.0ps
X258 X246-LSmitll_OR2T-OUT-X258-LSmitll_SPLITT-IN X258-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-INt X258-LSmitll_SPLITT-OUT-X265-LSmitll_DFFT-INt LSmitll_SPLITT

t1220 X259-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-INt 0 X259-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1221 X259-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt 0 X259-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN 0 z0=5 td=4.9ps
X259 X247-LSmitll_DFFT-OUT-X259-LSmitll_SPLITT-IN X259-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-INt X259-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt LSmitll_SPLITT

t1222 X260-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-INt 0 X260-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-IN 0 z0=5 td=8.7ps
t1223 X260-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-INt 0 X260-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-IN 0 z0=5 td=3.2ps
X260 X253-LSmitll_DFFT-OUT-X260-LSmitll_SPLITT-IN X260-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-INt X260-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-INt LSmitll_SPLITT

t1224 X261-LSmitll_DFFT-OUT-X275-LSmitll_SPLITT-INt 0 X261-LSmitll_DFFT-OUT-X275-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X261 X256-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-IN X456-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-IN X261-LSmitll_DFFT-OUT-X275-LSmitll_SPLITT-INt LSmitll_DFFT

t1225 X262-LSmitll_DFFT-OUT-X277-LSmitll_DFFT-INt 0 X262-LSmitll_DFFT-OUT-X277-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X262 X243-LSmitll_DFFT-OUT-X262-LSmitll_DFFT-IN X459-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-IN X262-LSmitll_DFFT-OUT-X277-LSmitll_DFFT-INt LSmitll_DFFT

t1226 X263-LSmitll_DFFT-OUT-X278-LSmitll_DFFT-INt 0 X263-LSmitll_DFFT-OUT-X278-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X263 X257-LSmitll_SPLITT-OUT-X263-LSmitll_DFFT-IN X551-LSmitll_SPLITT-OUT-X263-LSmitll_DFFT-IN X263-LSmitll_DFFT-OUT-X278-LSmitll_DFFT-INt LSmitll_DFFT

t1227 X264-LSmitll_DFFT-OUT-X279-LSmitll_DFFT-INt 0 X264-LSmitll_DFFT-OUT-X279-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X264 X245-LSmitll_DFFT-OUT-X264-LSmitll_DFFT-IN X348-LSmitll_SPLITT-OUT-X264-LSmitll_DFFT-IN X264-LSmitll_DFFT-OUT-X279-LSmitll_DFFT-INt LSmitll_DFFT

t1228 X265-LSmitll_DFFT-OUT-X280-LSmitll_OR2T-INt 0 X265-LSmitll_DFFT-OUT-X280-LSmitll_OR2T-IN 0 z0=5 td=2.4ps
X265 X258-LSmitll_SPLITT-OUT-X265-LSmitll_DFFT-IN X552-LSmitll_SPLITT-OUT-X265-LSmitll_DFFT-IN X265-LSmitll_DFFT-OUT-X280-LSmitll_OR2T-INt LSmitll_DFFT

t1229 X266-LSmitll_AND2T-OUT-X280-LSmitll_OR2T-INt 0 X266-LSmitll_AND2T-OUT-X280-LSmitll_OR2T-IN 0 z0=5 td=4.3ps
X266 X256-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN X259-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN X356-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN X266-LSmitll_AND2T-OUT-X280-LSmitll_OR2T-INt LSmitll_AND2T

t1230 X267-LSmitll_DFFT-OUT-X281-LSmitll_DFFT-INt 0 X267-LSmitll_DFFT-OUT-X281-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X267 X248-LSmitll_DFFT-OUT-X267-LSmitll_DFFT-IN X453-LSmitll_SPLITT-OUT-X267-LSmitll_DFFT-IN X267-LSmitll_DFFT-OUT-X281-LSmitll_DFFT-INt LSmitll_DFFT

t1231 X268-LSmitll_DFFT-OUT-X282-LSmitll_OR2T-INt 0 X268-LSmitll_DFFT-OUT-X282-LSmitll_OR2T-IN 0 z0=5 td=1.0ps
X268 X249-LSmitll_OR2T-OUT-X268-LSmitll_DFFT-IN X468-LSmitll_SPLITT-OUT-X268-LSmitll_DFFT-IN X268-LSmitll_DFFT-OUT-X282-LSmitll_OR2T-INt LSmitll_DFFT

t1232 X269-LSmitll_AND2T-OUT-X282-LSmitll_OR2T-INt 0 X269-LSmitll_AND2T-OUT-X282-LSmitll_OR2T-IN 0 z0=5 td=10.6ps
X269 X250-LSmitll_DFFT-OUT-X269-LSmitll_AND2T-IN X257-LSmitll_SPLITT-OUT-X269-LSmitll_AND2T-IN X351-LSmitll_SPLITT-OUT-X269-LSmitll_AND2T-IN X269-LSmitll_AND2T-OUT-X282-LSmitll_OR2T-INt LSmitll_AND2T

t1233 X270-LSmitll_DFFT-OUT-X283-LSmitll_DFFT-INt 0 X270-LSmitll_DFFT-OUT-X283-LSmitll_DFFT-IN 0 z0=5 td=6.6ps
X270 X251-LSmitll_DFFT-OUT-X270-LSmitll_DFFT-IN X456-LSmitll_SPLITT-OUT-X270-LSmitll_DFFT-IN X270-LSmitll_DFFT-OUT-X283-LSmitll_DFFT-INt LSmitll_DFFT

t1234 X271-LSmitll_DFFT-OUT-X284-LSmitll_OR2T-INt 0 X271-LSmitll_DFFT-OUT-X284-LSmitll_OR2T-IN 0 z0=5 td=4.6ps
X271 X252-LSmitll_OR2T-OUT-X271-LSmitll_DFFT-IN X394-LSmitll_SPLITT-OUT-X271-LSmitll_DFFT-IN X271-LSmitll_DFFT-OUT-X284-LSmitll_OR2T-INt LSmitll_DFFT

t1235 X272-LSmitll_AND2T-OUT-X284-LSmitll_OR2T-INt 0 X272-LSmitll_AND2T-OUT-X284-LSmitll_OR2T-IN 0 z0=5 td=12.5ps
X272 X258-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-IN X260-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-IN X369-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-IN X272-LSmitll_AND2T-OUT-X284-LSmitll_OR2T-INt LSmitll_AND2T

t1236 X273-LSmitll_AND2T-OUT-X285-LSmitll_AND2T-INt 0 X273-LSmitll_AND2T-OUT-X285-LSmitll_AND2T-IN 0 z0=5 td=10.9ps
X273 X259-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-IN X260-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-IN X553-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-IN X273-LSmitll_AND2T-OUT-X285-LSmitll_AND2T-INt LSmitll_AND2T

t1237 X274-LSmitll_DFFT-OUT-X286-LSmitll_DFFT-INt 0 X274-LSmitll_DFFT-OUT-X286-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X274 X254-LSmitll_AND2T-OUT-X274-LSmitll_DFFT-IN X467-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-IN X274-LSmitll_DFFT-OUT-X286-LSmitll_DFFT-INt LSmitll_DFFT

t1238 X275-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-INt 0 X275-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-IN 0 z0=5 td=8.5ps
t1239 X275-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-INt 0 X275-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-IN 0 z0=5 td=3.6ps
X275 X261-LSmitll_DFFT-OUT-X275-LSmitll_SPLITT-IN X275-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-INt X275-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-INt LSmitll_SPLITT

t1240 X276-LSmitll_DFFT-OUT-X288-LSmitll_XORT-INt 0 X276-LSmitll_DFFT-OUT-X288-LSmitll_XORT-IN 0 z0=5 td=2.6ps
X276 X275-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-IN X434-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-IN X276-LSmitll_DFFT-OUT-X288-LSmitll_XORT-INt LSmitll_DFFT

t1241 X277-LSmitll_DFFT-OUT-X288-LSmitll_XORT-INt 0 X277-LSmitll_DFFT-OUT-X288-LSmitll_XORT-IN 0 z0=5 td=1.0ps
X277 X262-LSmitll_DFFT-OUT-X277-LSmitll_DFFT-IN X454-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-IN X277-LSmitll_DFFT-OUT-X288-LSmitll_XORT-INt LSmitll_DFFT

t1242 X278-LSmitll_DFFT-OUT-X289-LSmitll_XORT-INt 0 X278-LSmitll_DFFT-OUT-X289-LSmitll_XORT-IN 0 z0=5 td=1.4ps
X278 X263-LSmitll_DFFT-OUT-X278-LSmitll_DFFT-IN X354-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-IN X278-LSmitll_DFFT-OUT-X289-LSmitll_XORT-INt LSmitll_DFFT

t1243 X279-LSmitll_DFFT-OUT-X289-LSmitll_XORT-INt 0 X279-LSmitll_DFFT-OUT-X289-LSmitll_XORT-IN 0 z0=5 td=2.4ps
X279 X264-LSmitll_DFFT-OUT-X279-LSmitll_DFFT-IN X349-LSmitll_SPLITT-OUT-X279-LSmitll_DFFT-IN X279-LSmitll_DFFT-OUT-X289-LSmitll_XORT-INt LSmitll_DFFT

t1244 X280-LSmitll_OR2T-OUT-X290-LSmitll_XORT-INt 0 X280-LSmitll_OR2T-OUT-X290-LSmitll_XORT-IN 0 z0=5 td=8.1ps
X280 X265-LSmitll_DFFT-OUT-X280-LSmitll_OR2T-IN X266-LSmitll_AND2T-OUT-X280-LSmitll_OR2T-IN X428-LSmitll_SPLITT-OUT-X280-LSmitll_OR2T-IN X280-LSmitll_OR2T-OUT-X290-LSmitll_XORT-INt LSmitll_OR2T

t1245 X281-LSmitll_DFFT-OUT-X290-LSmitll_XORT-INt 0 X281-LSmitll_DFFT-OUT-X290-LSmitll_XORT-IN 0 z0=5 td=3.5ps
X281 X267-LSmitll_DFFT-OUT-X281-LSmitll_DFFT-IN X554-LSmitll_SPLITT-OUT-X281-LSmitll_DFFT-IN X281-LSmitll_DFFT-OUT-X290-LSmitll_XORT-INt LSmitll_DFFT

t1246 X282-LSmitll_OR2T-OUT-X287-LSmitll_SPLITT-INt 0 X282-LSmitll_OR2T-OUT-X287-LSmitll_SPLITT-IN 0 z0=5 td=12.1ps
X282 X268-LSmitll_DFFT-OUT-X282-LSmitll_OR2T-IN X269-LSmitll_AND2T-OUT-X282-LSmitll_OR2T-IN X431-LSmitll_SPLITT-OUT-X282-LSmitll_OR2T-IN X282-LSmitll_OR2T-OUT-X287-LSmitll_SPLITT-INt LSmitll_OR2T

t1247 X283-LSmitll_DFFT-OUT-X291-LSmitll_XORT-INt 0 X283-LSmitll_DFFT-OUT-X291-LSmitll_XORT-IN 0 z0=5 td=2.4ps
X283 X270-LSmitll_DFFT-OUT-X283-LSmitll_DFFT-IN X459-LSmitll_SPLITT-OUT-X283-LSmitll_DFFT-IN X283-LSmitll_DFFT-OUT-X291-LSmitll_XORT-INt LSmitll_DFFT

t1248 X284-LSmitll_OR2T-OUT-X292-LSmitll_OR2T-INt 0 X284-LSmitll_OR2T-OUT-X292-LSmitll_OR2T-IN 0 z0=5 td=2.6ps
X284 X271-LSmitll_DFFT-OUT-X284-LSmitll_OR2T-IN X272-LSmitll_AND2T-OUT-X284-LSmitll_OR2T-IN X356-LSmitll_SPLITT-OUT-X284-LSmitll_OR2T-IN X284-LSmitll_OR2T-OUT-X292-LSmitll_OR2T-INt LSmitll_OR2T

t1249 X285-LSmitll_AND2T-OUT-X292-LSmitll_OR2T-INt 0 X285-LSmitll_AND2T-OUT-X292-LSmitll_OR2T-IN 0 z0=5 td=5.4ps
X285 X273-LSmitll_AND2T-OUT-X285-LSmitll_AND2T-IN X275-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-IN X431-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-IN X285-LSmitll_AND2T-OUT-X292-LSmitll_OR2T-INt LSmitll_AND2T

t1250 X286-LSmitll_DFFT-OUT-X294-LSmitll_DFFT-INt 0 X286-LSmitll_DFFT-OUT-X294-LSmitll_DFFT-IN 0 z0=5 td=8.5ps
X286 X274-LSmitll_DFFT-OUT-X286-LSmitll_DFFT-IN X555-LSmitll_SPLITT-OUT-X286-LSmitll_DFFT-IN X286-LSmitll_DFFT-OUT-X294-LSmitll_DFFT-INt LSmitll_DFFT

t1251 X287-LSmitll_SPLITT-OUT-X293-LSmitll_DFFT-INt 0 X287-LSmitll_SPLITT-OUT-X293-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t1252 X287-LSmitll_SPLITT-OUT-X291-LSmitll_XORT-INt 0 X287-LSmitll_SPLITT-OUT-X291-LSmitll_XORT-IN 0 z0=5 td=4.1ps
X287 X282-LSmitll_OR2T-OUT-X287-LSmitll_SPLITT-IN X287-LSmitll_SPLITT-OUT-X293-LSmitll_DFFT-INt X287-LSmitll_SPLITT-OUT-X291-LSmitll_XORT-INt LSmitll_SPLITT

t1253 X288-LSmitll_XORT-OUT-X301-LSmitll_DFFT-INt 0 X288-LSmitll_XORT-OUT-X301-LSmitll_DFFT-IN 0 z0=5 td=7.9ps
X288 X276-LSmitll_DFFT-OUT-X288-LSmitll_XORT-IN X277-LSmitll_DFFT-OUT-X288-LSmitll_XORT-IN X453-LSmitll_SPLITT-OUT-X288-LSmitll_XORT-IN X288-LSmitll_XORT-OUT-X301-LSmitll_DFFT-INt LSmitll_XORT

t1254 X289-LSmitll_XORT-OUT-X300-LSmitll_DFFT-INt 0 X289-LSmitll_XORT-OUT-X300-LSmitll_DFFT-IN 0 z0=5 td=12.4ps
X289 X278-LSmitll_DFFT-OUT-X289-LSmitll_XORT-IN X279-LSmitll_DFFT-OUT-X289-LSmitll_XORT-IN X354-LSmitll_SPLITT-OUT-X289-LSmitll_XORT-IN X289-LSmitll_XORT-OUT-X300-LSmitll_DFFT-INt LSmitll_XORT

t1255 X290-LSmitll_XORT-OUT-X299-LSmitll_DFFT-INt 0 X290-LSmitll_XORT-OUT-X299-LSmitll_DFFT-IN 0 z0=5 td=7.1ps
X290 X280-LSmitll_OR2T-OUT-X290-LSmitll_XORT-IN X281-LSmitll_DFFT-OUT-X290-LSmitll_XORT-IN X556-LSmitll_SPLITT-OUT-X290-LSmitll_XORT-IN X290-LSmitll_XORT-OUT-X299-LSmitll_DFFT-INt LSmitll_XORT

t1256 X291-LSmitll_XORT-OUT-X295-LSmitll_SPLITT-INt 0 X291-LSmitll_XORT-OUT-X295-LSmitll_SPLITT-IN 0 z0=5 td=6.3ps
X291 X283-LSmitll_DFFT-OUT-X291-LSmitll_XORT-IN X287-LSmitll_SPLITT-OUT-X291-LSmitll_XORT-IN X461-LSmitll_SPLITT-OUT-X291-LSmitll_XORT-IN X291-LSmitll_XORT-OUT-X295-LSmitll_SPLITT-INt LSmitll_XORT

t1257 X292-LSmitll_OR2T-OUT-X296-LSmitll_XORT-INt 0 X292-LSmitll_OR2T-OUT-X296-LSmitll_XORT-IN 0 z0=5 td=9.2ps
X292 X284-LSmitll_OR2T-OUT-X292-LSmitll_OR2T-IN X285-LSmitll_AND2T-OUT-X292-LSmitll_OR2T-IN X557-LSmitll_SPLITT-OUT-X292-LSmitll_OR2T-IN X292-LSmitll_OR2T-OUT-X296-LSmitll_XORT-INt LSmitll_OR2T

t1258 X293-LSmitll_DFFT-OUT-X296-LSmitll_XORT-INt 0 X293-LSmitll_DFFT-OUT-X296-LSmitll_XORT-IN 0 z0=5 td=2.6ps
X293 X287-LSmitll_SPLITT-OUT-X293-LSmitll_DFFT-IN X558-LSmitll_SPLITT-OUT-X293-LSmitll_DFFT-IN X293-LSmitll_DFFT-OUT-X296-LSmitll_XORT-INt LSmitll_DFFT

t1259 X294-LSmitll_DFFT-OUT-X302-LSmitll_DFFT-INt 0 X294-LSmitll_DFFT-OUT-X302-LSmitll_DFFT-IN 0 z0=5 td=3.7ps
X294 X286-LSmitll_DFFT-OUT-X294-LSmitll_DFFT-IN X492-LSmitll_SPLITT-OUT-X294-LSmitll_DFFT-IN X294-LSmitll_DFFT-OUT-X302-LSmitll_DFFT-INt LSmitll_DFFT

t1260 X295-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-INt 0 X295-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-IN 0 z0=5 td=3.3ps
t1261 X295-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-INt 0 X295-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
X295 X291-LSmitll_XORT-OUT-X295-LSmitll_SPLITT-IN X295-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-INt X295-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-INt LSmitll_SPLITT

t1262 X296-LSmitll_XORT-OUT-X307-LSmitll_DFFT-INt 0 X296-LSmitll_XORT-OUT-X307-LSmitll_DFFT-IN 0 z0=5 td=4.1ps
X296 X292-LSmitll_OR2T-OUT-X296-LSmitll_XORT-IN X293-LSmitll_DFFT-OUT-X296-LSmitll_XORT-IN X461-LSmitll_SPLITT-OUT-X296-LSmitll_XORT-IN X296-LSmitll_XORT-OUT-X307-LSmitll_DFFT-INt LSmitll_XORT

t1263 X297-LSmitll_DFFT-OUT-X309-LSmitll_DFFT-INt 0 X297-LSmitll_DFFT-OUT-X309-LSmitll_DFFT-IN 0 z0=5 td=5.6ps
X297 X295-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-IN X559-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-IN X297-LSmitll_DFFT-OUT-X309-LSmitll_DFFT-INt LSmitll_DFFT

t1264 X298-LSmitll_DFFT-OUT-X303-LSmitll_DFFT-INt 0 X298-LSmitll_DFFT-OUT-X303-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X298 X295-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-IN X449-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-IN X298-LSmitll_DFFT-OUT-X303-LSmitll_DFFT-INt LSmitll_DFFT

t1265 X299-LSmitll_DFFT-OUT-X304-LSmitll_DFFT-INt 0 X299-LSmitll_DFFT-OUT-X304-LSmitll_DFFT-IN 0 z0=5 td=6.1ps
X299 X290-LSmitll_XORT-OUT-X299-LSmitll_DFFT-IN X560-LSmitll_SPLITT-OUT-X299-LSmitll_DFFT-IN X299-LSmitll_DFFT-OUT-X304-LSmitll_DFFT-INt LSmitll_DFFT

t1266 X300-LSmitll_DFFT-OUT-X305-LSmitll_DFFT-INt 0 X300-LSmitll_DFFT-OUT-X305-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X300 X289-LSmitll_XORT-OUT-X300-LSmitll_DFFT-IN X316-LSmitll_SPLITT-OUT-X300-LSmitll_DFFT-IN X300-LSmitll_DFFT-OUT-X305-LSmitll_DFFT-INt LSmitll_DFFT

t1267 X301-LSmitll_DFFT-OUT-X306-LSmitll_DFFT-INt 0 X301-LSmitll_DFFT-OUT-X306-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X301 X288-LSmitll_XORT-OUT-X301-LSmitll_DFFT-IN X336-LSmitll_SPLITT-OUT-X301-LSmitll_DFFT-IN X301-LSmitll_DFFT-OUT-X306-LSmitll_DFFT-INt LSmitll_DFFT

t1268 X302-LSmitll_DFFT-OUT-X308-LSmitll_DFFT-INt 0 X302-LSmitll_DFFT-OUT-X308-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X302 X294-LSmitll_DFFT-OUT-X302-LSmitll_DFFT-IN X561-LSmitll_SPLITT-OUT-X302-LSmitll_DFFT-IN X302-LSmitll_DFFT-OUT-X308-LSmitll_DFFT-INt LSmitll_DFFT

t1269 X303-LSmitll_DFFT-OUT-X58-LSmitll_AND2T-INt 0 X303-LSmitll_DFFT-OUT-X58-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
X303 X298-LSmitll_DFFT-OUT-X303-LSmitll_DFFT-IN X447-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-IN X303-LSmitll_DFFT-OUT-X58-LSmitll_AND2T-INt LSmitll_DFFT

t1270 X304-LSmitll_DFFT-OUT-X60-LSmitll_AND2T-INt 0 X304-LSmitll_DFFT-OUT-X60-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
X304 X299-LSmitll_DFFT-OUT-X304-LSmitll_DFFT-IN X562-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-IN X304-LSmitll_DFFT-OUT-X60-LSmitll_AND2T-INt LSmitll_DFFT

t1271 X305-LSmitll_DFFT-OUT-X62-LSmitll_AND2T-INt 0 X305-LSmitll_DFFT-OUT-X62-LSmitll_AND2T-IN 0 z0=5 td=11.7ps
X305 X300-LSmitll_DFFT-OUT-X305-LSmitll_DFFT-IN X316-LSmitll_SPLITT-OUT-X305-LSmitll_DFFT-IN X305-LSmitll_DFFT-OUT-X62-LSmitll_AND2T-INt LSmitll_DFFT

t1272 X306-LSmitll_DFFT-OUT-X64-LSmitll_AND2T-INt 0 X306-LSmitll_DFFT-OUT-X64-LSmitll_AND2T-IN 0 z0=5 td=5.0ps
X306 X301-LSmitll_DFFT-OUT-X306-LSmitll_DFFT-IN X337-LSmitll_SPLITT-OUT-X306-LSmitll_DFFT-IN X306-LSmitll_DFFT-OUT-X64-LSmitll_AND2T-INt LSmitll_DFFT

t1273 X307-LSmitll_DFFT-OUT-X110-LSmitll_AND2T-INt 0 X307-LSmitll_DFFT-OUT-X110-LSmitll_AND2T-IN 0 z0=5 td=3.3ps
X307 X296-LSmitll_XORT-OUT-X307-LSmitll_DFFT-IN X563-LSmitll_SPLITT-OUT-X307-LSmitll_DFFT-IN X307-LSmitll_DFFT-OUT-X110-LSmitll_AND2T-INt LSmitll_DFFT

t1274 X308-LSmitll_DFFT-OUT-X113-LSmitll_AND2T-INt 0 X308-LSmitll_DFFT-OUT-X113-LSmitll_AND2T-IN 0 z0=5 td=5.8ps
X308 X302-LSmitll_DFFT-OUT-X308-LSmitll_DFFT-IN X495-LSmitll_SPLITT-OUT-X308-LSmitll_DFFT-IN X308-LSmitll_DFFT-OUT-X113-LSmitll_AND2T-INt LSmitll_DFFT

t1275 X309-LSmitll_DFFT-OUT-X116-LSmitll_AND2T-INt 0 X309-LSmitll_DFFT-OUT-X116-LSmitll_AND2T-IN 0 z0=5 td=2.7ps
X309 X297-LSmitll_DFFT-OUT-X309-LSmitll_DFFT-IN X424-LSmitll_SPLITT-OUT-X309-LSmitll_DFFT-IN X309-LSmitll_DFFT-OUT-X116-LSmitll_AND2T-INt LSmitll_DFFT

t1276 X310-LSmitll_SPLITT-OUT-X61-LSmitll_AND2T-INt 0 X310-LSmitll_SPLITT-OUT-X61-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
t1277 X310-LSmitll_SPLITT-OUT-X75-LSmitll_OR2T-INt 0 X310-LSmitll_SPLITT-OUT-X75-LSmitll_OR2T-IN 0 z0=5 td=0.5ps
X310 X312-LSmitll_SPLITT-OUT-X310-LSmitll_SPLITT-IN X310-LSmitll_SPLITT-OUT-X61-LSmitll_AND2T-INt X310-LSmitll_SPLITT-OUT-X75-LSmitll_OR2T-INt LSmitll_SPLITT

t1278 X311-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-INt 0 X311-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
t1279 X311-LSmitll_SPLITT-OUT-X62-LSmitll_AND2T-INt 0 X311-LSmitll_SPLITT-OUT-X62-LSmitll_AND2T-IN 0 z0=5 td=0.8ps
X311 X312-LSmitll_SPLITT-OUT-X311-LSmitll_SPLITT-IN X311-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-INt X311-LSmitll_SPLITT-OUT-X62-LSmitll_AND2T-INt LSmitll_SPLITT

t1280 X312-LSmitll_SPLITT-OUT-X310-LSmitll_SPLITT-INt 0 X312-LSmitll_SPLITT-OUT-X310-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1281 X312-LSmitll_SPLITT-OUT-X311-LSmitll_SPLITT-INt 0 X312-LSmitll_SPLITT-OUT-X311-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X312 X315-LSmitll_SPLITT-OUT-X312-LSmitll_SPLITT-IN X312-LSmitll_SPLITT-OUT-X310-LSmitll_SPLITT-INt X312-LSmitll_SPLITT-OUT-X311-LSmitll_SPLITT-INt LSmitll_SPLITT

t1282 X313-LSmitll_SPLITT-OUT-X37-LSmitll_DFFT-INt 0 X313-LSmitll_SPLITT-OUT-X37-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
t1283 X313-LSmitll_SPLITT-OUT-X38-LSmitll_DFFT-INt 0 X313-LSmitll_SPLITT-OUT-X38-LSmitll_DFFT-IN 0 z0=5 td=4.0ps
X313 X314-LSmitll_SPLITT-OUT-X313-LSmitll_SPLITT-IN X313-LSmitll_SPLITT-OUT-X37-LSmitll_DFFT-INt X313-LSmitll_SPLITT-OUT-X38-LSmitll_DFFT-INt LSmitll_SPLITT

t1284 X314-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-INt 0 X314-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1285 X314-LSmitll_SPLITT-OUT-X313-LSmitll_SPLITT-INt 0 X314-LSmitll_SPLITT-OUT-X313-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X314 X315-LSmitll_SPLITT-OUT-X314-LSmitll_SPLITT-IN X314-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-INt X314-LSmitll_SPLITT-OUT-X313-LSmitll_SPLITT-INt LSmitll_SPLITT

t1286 X315-LSmitll_SPLITT-OUT-X312-LSmitll_SPLITT-INt 0 X315-LSmitll_SPLITT-OUT-X312-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1287 X315-LSmitll_SPLITT-OUT-X314-LSmitll_SPLITT-INt 0 X315-LSmitll_SPLITT-OUT-X314-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X315 X322-LSmitll_SPLITT-OUT-X315-LSmitll_SPLITT-IN X315-LSmitll_SPLITT-OUT-X312-LSmitll_SPLITT-INt X315-LSmitll_SPLITT-OUT-X314-LSmitll_SPLITT-INt LSmitll_SPLITT

t1288 X316-LSmitll_SPLITT-OUT-X300-LSmitll_DFFT-INt 0 X316-LSmitll_SPLITT-OUT-X300-LSmitll_DFFT-IN 0 z0=5 td=1.7ps
t1289 X316-LSmitll_SPLITT-OUT-X305-LSmitll_DFFT-INt 0 X316-LSmitll_SPLITT-OUT-X305-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
X316 X318-LSmitll_SPLITT-OUT-X316-LSmitll_SPLITT-IN X316-LSmitll_SPLITT-OUT-X300-LSmitll_DFFT-INt X316-LSmitll_SPLITT-OUT-X305-LSmitll_DFFT-INt LSmitll_SPLITT

t1290 X317-LSmitll_SPLITT-OUT-X27-LSmitll_NOTT-INt 0 X317-LSmitll_SPLITT-OUT-X27-LSmitll_NOTT-IN 0 z0=5 td=2.3ps
t1291 X317-LSmitll_SPLITT-OUT-X36-LSmitll_DFFT-INt 0 X317-LSmitll_SPLITT-OUT-X36-LSmitll_DFFT-IN 0 z0=5 td=2.4ps
X317 X318-LSmitll_SPLITT-OUT-X317-LSmitll_SPLITT-IN X317-LSmitll_SPLITT-OUT-X27-LSmitll_NOTT-INt X317-LSmitll_SPLITT-OUT-X36-LSmitll_DFFT-INt LSmitll_SPLITT

t1292 X318-LSmitll_SPLITT-OUT-X316-LSmitll_SPLITT-INt 0 X318-LSmitll_SPLITT-OUT-X316-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1293 X318-LSmitll_SPLITT-OUT-X317-LSmitll_SPLITT-INt 0 X318-LSmitll_SPLITT-OUT-X317-LSmitll_SPLITT-IN 0 z0=5 td=0.5ps
X318 X321-LSmitll_SPLITT-OUT-X318-LSmitll_SPLITT-IN X318-LSmitll_SPLITT-OUT-X316-LSmitll_SPLITT-INt X318-LSmitll_SPLITT-OUT-X317-LSmitll_SPLITT-INt LSmitll_SPLITT

t1294 X319-LSmitll_SPLITT-OUT-X97-LSmitll_NDROT-INt 0 X319-LSmitll_SPLITT-OUT-X97-LSmitll_NDROT-IN 0 z0=5 td=3.6ps
t1295 X319-LSmitll_SPLITT-OUT-X103-LSmitll_NDROT-INt 0 X319-LSmitll_SPLITT-OUT-X103-LSmitll_NDROT-IN 0 z0=5 td=0.8ps
X319 X320-LSmitll_SPLITT-OUT-X319-LSmitll_SPLITT-IN X319-LSmitll_SPLITT-OUT-X97-LSmitll_NDROT-INt X319-LSmitll_SPLITT-OUT-X103-LSmitll_NDROT-INt LSmitll_SPLITT

t1296 X320-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-INt 0 X320-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1297 X320-LSmitll_SPLITT-OUT-X319-LSmitll_SPLITT-INt 0 X320-LSmitll_SPLITT-OUT-X319-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X320 X321-LSmitll_SPLITT-OUT-X320-LSmitll_SPLITT-IN X320-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-INt X320-LSmitll_SPLITT-OUT-X319-LSmitll_SPLITT-INt LSmitll_SPLITT

t1298 X321-LSmitll_SPLITT-OUT-X318-LSmitll_SPLITT-INt 0 X321-LSmitll_SPLITT-OUT-X318-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1299 X321-LSmitll_SPLITT-OUT-X320-LSmitll_SPLITT-INt 0 X321-LSmitll_SPLITT-OUT-X320-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X321 X322-LSmitll_SPLITT-OUT-X321-LSmitll_SPLITT-IN X321-LSmitll_SPLITT-OUT-X318-LSmitll_SPLITT-INt X321-LSmitll_SPLITT-OUT-X320-LSmitll_SPLITT-INt LSmitll_SPLITT

t1300 X322-LSmitll_SPLITT-OUT-X315-LSmitll_SPLITT-INt 0 X322-LSmitll_SPLITT-OUT-X315-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1301 X322-LSmitll_SPLITT-OUT-X321-LSmitll_SPLITT-INt 0 X322-LSmitll_SPLITT-OUT-X321-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
X322 X335-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-IN X322-LSmitll_SPLITT-OUT-X315-LSmitll_SPLITT-INt X322-LSmitll_SPLITT-OUT-X321-LSmitll_SPLITT-INt LSmitll_SPLITT

t1302 X323-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-INt 0 X323-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1303 X323-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-INt 0 X323-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
X323 X325-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-IN X323-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-INt X323-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-INt LSmitll_SPLITT

t1304 X324-LSmitll_SPLITT-OUT-X100-LSmitll_NDROT-INt 0 X324-LSmitll_SPLITT-OUT-X100-LSmitll_NDROT-IN 0 z0=5 td=3.0ps
t1305 X324-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt 0 X324-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
X324 X325-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-IN X324-LSmitll_SPLITT-OUT-X100-LSmitll_NDROT-INt X324-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt LSmitll_SPLITT

t1306 X325-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-INt 0 X325-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
t1307 X325-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-INt 0 X325-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X325 X328-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-IN X325-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-INt X325-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-INt LSmitll_SPLITT

t1308 X326-LSmitll_SPLITT-OUT-X198-LSmitll_DFFT-INt 0 X326-LSmitll_SPLITT-OUT-X198-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
t1309 X326-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-INt 0 X326-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-IN 0 z0=5 td=2.0ps
X326 X327-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-IN X326-LSmitll_SPLITT-OUT-X198-LSmitll_DFFT-INt X326-LSmitll_SPLITT-OUT-X242-LSmitll_DFFT-INt LSmitll_SPLITT

t1310 X327-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-INt 0 X327-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1311 X327-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-INt 0 X327-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X327 X328-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-IN X327-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-INt X327-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-INt LSmitll_SPLITT

t1312 X328-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-INt 0 X328-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1313 X328-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-INt 0 X328-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X328 X334-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-IN X328-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-INt X328-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-INt LSmitll_SPLITT

t1314 X329-LSmitll_SPLITT-OUT-X229-LSmitll_DFFT-INt 0 X329-LSmitll_SPLITT-OUT-X229-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
t1315 X329-LSmitll_SPLITT-OUT-X255-LSmitll_DFFT-INt 0 X329-LSmitll_SPLITT-OUT-X255-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
X329 X330-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-IN X329-LSmitll_SPLITT-OUT-X229-LSmitll_DFFT-INt X329-LSmitll_SPLITT-OUT-X255-LSmitll_DFFT-INt LSmitll_SPLITT

t1316 X330-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-INt 0 X330-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1317 X330-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-INt 0 X330-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
X330 X333-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-IN X330-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-INt X330-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-INt LSmitll_SPLITT

t1318 X331-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-INt 0 X331-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-IN 0 z0=5 td=3.2ps
t1319 X331-LSmitll_SPLITT-OUT-X246-LSmitll_OR2T-INt 0 X331-LSmitll_SPLITT-OUT-X246-LSmitll_OR2T-IN 0 z0=5 td=2.8ps
X331 X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-IN X331-LSmitll_SPLITT-OUT-X227-LSmitll_AND2T-INt X331-LSmitll_SPLITT-OUT-X246-LSmitll_OR2T-INt LSmitll_SPLITT

t1320 X332-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-INt 0 X332-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-IN 0 z0=5 td=4.0ps
t1321 X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-INt 0 X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X332 X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-IN X332-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-INt X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-INt LSmitll_SPLITT

t1322 X333-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-INt 0 X333-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1323 X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-INt 0 X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X333 X334-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-IN X333-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-INt X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-INt LSmitll_SPLITT

t1324 X334-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-INt 0 X334-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1325 X334-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-INt 0 X334-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X334 X335-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-IN X334-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-INt X334-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-INt LSmitll_SPLITT

t1326 X335-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-INt 0 X335-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1327 X335-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-INt 0 X335-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X335 X361-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-IN X335-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-INt X335-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-INt LSmitll_SPLITT

t1328 X336-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-INt 0 X336-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-IN 0 z0=5 td=4.0ps
t1329 X336-LSmitll_SPLITT-OUT-X301-LSmitll_DFFT-INt 0 X336-LSmitll_SPLITT-OUT-X301-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X336 X338-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-IN X336-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-INt X336-LSmitll_SPLITT-OUT-X301-LSmitll_DFFT-INt LSmitll_SPLITT

t1330 X337-LSmitll_SPLITT-OUT-X29-LSmitll_NOTT-INt 0 X337-LSmitll_SPLITT-OUT-X29-LSmitll_NOTT-IN 0 z0=5 td=2.5ps
t1331 X337-LSmitll_SPLITT-OUT-X306-LSmitll_DFFT-INt 0 X337-LSmitll_SPLITT-OUT-X306-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
X337 X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-IN X337-LSmitll_SPLITT-OUT-X29-LSmitll_NOTT-INt X337-LSmitll_SPLITT-OUT-X306-LSmitll_DFFT-INt LSmitll_SPLITT

t1332 X338-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-INt 0 X338-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1333 X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-INt 0 X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X338 X341-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-IN X338-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-INt X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-INt LSmitll_SPLITT

t1334 X339-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-INt 0 X339-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-IN 0 z0=5 td=2.4ps
t1335 X339-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt 0 X339-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN 0 z0=5 td=1.3ps
X339 X340-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-IN X339-LSmitll_SPLITT-OUT-X79-LSmitll_DFFT-INt X339-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt LSmitll_SPLITT

t1336 X340-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-INt 0 X340-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1337 X340-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-INt 0 X340-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X340 X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-IN X340-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-INt X340-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-INt LSmitll_SPLITT

t1338 X341-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-INt 0 X341-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1339 X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-INt 0 X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
X341 X347-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-IN X341-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-INt X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-INt LSmitll_SPLITT

t1340 X342-LSmitll_SPLITT-OUT-X6-LSmitll_DFFT-INt 0 X342-LSmitll_SPLITT-OUT-X6-LSmitll_DFFT-IN 0 z0=5 td=2.5ps
t1341 X342-LSmitll_SPLITT-OUT-X64-LSmitll_AND2T-INt 0 X342-LSmitll_SPLITT-OUT-X64-LSmitll_AND2T-IN 0 z0=5 td=0.7ps
X342 X343-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-IN X342-LSmitll_SPLITT-OUT-X6-LSmitll_DFFT-INt X342-LSmitll_SPLITT-OUT-X64-LSmitll_AND2T-INt LSmitll_SPLITT

t1342 X343-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-INt 0 X343-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t1343 X343-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-INt 0 X343-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X343 X346-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-IN X343-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-INt X343-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-INt LSmitll_SPLITT

t1344 X344-LSmitll_SPLITT-OUT-X35-LSmitll_DFFT-INt 0 X344-LSmitll_SPLITT-OUT-X35-LSmitll_DFFT-IN 0 z0=5 td=5.7ps
t1345 X344-LSmitll_SPLITT-OUT-X40-LSmitll_DFFT-INt 0 X344-LSmitll_SPLITT-OUT-X40-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X344 X345-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-IN X344-LSmitll_SPLITT-OUT-X35-LSmitll_DFFT-INt X344-LSmitll_SPLITT-OUT-X40-LSmitll_DFFT-INt LSmitll_SPLITT

t1346 X345-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-INt 0 X345-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1347 X345-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-INt 0 X345-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X345 X346-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-IN X345-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-INt X345-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-INt LSmitll_SPLITT

t1348 X346-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-INt 0 X346-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1349 X346-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-INt 0 X346-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X346 X347-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-IN X346-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-INt X346-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-INt LSmitll_SPLITT

t1350 X347-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-INt 0 X347-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1351 X347-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-INt 0 X347-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X347 X360-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-IN X347-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-INt X347-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-INt LSmitll_SPLITT

t1352 X348-LSmitll_SPLITT-OUT-X245-LSmitll_DFFT-INt 0 X348-LSmitll_SPLITT-OUT-X245-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1353 X348-LSmitll_SPLITT-OUT-X264-LSmitll_DFFT-INt 0 X348-LSmitll_SPLITT-OUT-X264-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
X348 X350-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-IN X348-LSmitll_SPLITT-OUT-X245-LSmitll_DFFT-INt X348-LSmitll_SPLITT-OUT-X264-LSmitll_DFFT-INt LSmitll_SPLITT

t1354 X349-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-INt 0 X349-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
t1355 X349-LSmitll_SPLITT-OUT-X279-LSmitll_DFFT-INt 0 X349-LSmitll_SPLITT-OUT-X279-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
X349 X350-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-IN X349-LSmitll_SPLITT-OUT-X226-LSmitll_DFFT-INt X349-LSmitll_SPLITT-OUT-X279-LSmitll_DFFT-INt LSmitll_SPLITT

t1356 X350-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-INt 0 X350-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1357 X350-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-INt 0 X350-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X350 X353-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-IN X350-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-INt X350-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-INt LSmitll_SPLITT

t1358 X351-LSmitll_SPLITT-OUT-X247-LSmitll_DFFT-INt 0 X351-LSmitll_SPLITT-OUT-X247-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
t1359 X351-LSmitll_SPLITT-OUT-X269-LSmitll_AND2T-INt 0 X351-LSmitll_SPLITT-OUT-X269-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
X351 X352-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-IN X351-LSmitll_SPLITT-OUT-X247-LSmitll_DFFT-INt X351-LSmitll_SPLITT-OUT-X269-LSmitll_AND2T-INt LSmitll_SPLITT

t1360 X352-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-INt 0 X352-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1361 X352-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-INt 0 X352-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X352 X353-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-IN X352-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-INt X352-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-INt LSmitll_SPLITT

t1362 X353-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-INt 0 X353-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1363 X353-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-INt 0 X353-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
X353 X359-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-IN X353-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-INt X353-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-INt LSmitll_SPLITT

t1364 X354-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-INt 0 X354-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
t1365 X354-LSmitll_SPLITT-OUT-X289-LSmitll_XORT-INt 0 X354-LSmitll_SPLITT-OUT-X289-LSmitll_XORT-IN 0 z0=5 td=1.5ps
X354 X355-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-IN X354-LSmitll_SPLITT-OUT-X278-LSmitll_DFFT-INt X354-LSmitll_SPLITT-OUT-X289-LSmitll_XORT-INt LSmitll_SPLITT

t1366 X355-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-INt 0 X355-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1367 X355-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-INt 0 X355-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X355 X358-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-IN X355-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-INt X355-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-INt LSmitll_SPLITT

t1368 X356-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt 0 X356-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN 0 z0=5 td=0.5ps
t1369 X356-LSmitll_SPLITT-OUT-X284-LSmitll_OR2T-INt 0 X356-LSmitll_SPLITT-OUT-X284-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X356 X357-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-IN X356-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt X356-LSmitll_SPLITT-OUT-X284-LSmitll_OR2T-INt LSmitll_SPLITT

t1370 X357-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-INt 0 X357-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1371 X357-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-INt 0 X357-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X357 X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-IN X357-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-INt X357-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-INt LSmitll_SPLITT

t1372 X358-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-INt 0 X358-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1373 X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-INt 0 X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X358 X359-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-IN X358-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-INt X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-INt LSmitll_SPLITT

t1374 X359-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-INt 0 X359-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1375 X359-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-INt 0 X359-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X359 X360-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-IN X359-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-INt X359-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-INt LSmitll_SPLITT

t1376 X360-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-INt 0 X360-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-IN 0 z0=5 td=3.2ps
t1377 X360-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-INt 0 X360-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-IN 0 z0=5 td=4.0ps
X360 X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-IN X360-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-INt X360-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-INt LSmitll_SPLITT

t1378 X361-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-INt 0 X361-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-IN 0 z0=5 td=7.1ps
t1379 X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-INt 0 X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-IN 0 z0=5 td=5.5ps
X361 X414-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-IN X361-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-INt X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-INt LSmitll_SPLITT

t1380 X362-LSmitll_SPLITT-OUT-X19-LSmitll_DFFT-INt 0 X362-LSmitll_SPLITT-OUT-X19-LSmitll_DFFT-IN 0 z0=5 td=4.1ps
t1381 X362-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-INt 0 X362-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-IN 0 z0=5 td=1.7ps
X362 X364-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-IN X362-LSmitll_SPLITT-OUT-X19-LSmitll_DFFT-INt X362-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-INt LSmitll_SPLITT

t1382 X363-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-INt 0 X363-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
t1383 X363-LSmitll_SPLITT-OUT-X199-LSmitll_DFFT-INt 0 X363-LSmitll_SPLITT-OUT-X199-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
X363 X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-IN X363-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-INt X363-LSmitll_SPLITT-OUT-X199-LSmitll_DFFT-INt LSmitll_SPLITT

t1384 X364-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-INt 0 X364-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
t1385 X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-INt 0 X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X364 X367-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-IN X364-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-INt X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-INt LSmitll_SPLITT

t1386 X365-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-INt 0 X365-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t1387 X365-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt 0 X365-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN 0 z0=5 td=1.4ps
X365 X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-IN X365-LSmitll_SPLITT-OUT-X201-LSmitll_DFFT-INt X365-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt LSmitll_SPLITT

t1388 X366-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-INt 0 X366-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1389 X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-INt 0 X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X366 X367-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-IN X366-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-INt X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-INt LSmitll_SPLITT

t1390 X367-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-INt 0 X367-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1391 X367-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-INt 0 X367-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X367 X374-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-IN X367-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-INt X367-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-INt LSmitll_SPLITT

t1392 X368-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-INt 0 X368-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-IN 0 z0=5 td=2.6ps
t1393 X368-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-INt 0 X368-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
X368 X370-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-IN X368-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-INt X368-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-INt LSmitll_SPLITT

t1394 X369-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-INt 0 X369-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-IN 0 z0=5 td=10.7ps
t1395 X369-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-INt 0 X369-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
X369 X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-IN X369-LSmitll_SPLITT-OUT-X241-LSmitll_AND2T-INt X369-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-INt LSmitll_SPLITT

t1396 X370-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-INt 0 X370-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1397 X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-INt 0 X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X370 X373-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-IN X370-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-INt X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-INt LSmitll_SPLITT

t1398 X371-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-INt 0 X371-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
t1399 X371-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-INt 0 X371-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-IN 0 z0=5 td=3.1ps
X371 X372-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-IN X371-LSmitll_SPLITT-OUT-X182-LSmitll_AND2T-INt X371-LSmitll_SPLITT-OUT-X186-LSmitll_AND2T-INt LSmitll_SPLITT

t1400 X372-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-INt 0 X372-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1401 X372-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-INt 0 X372-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X372 X373-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-IN X372-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-INt X372-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-INt LSmitll_SPLITT

t1402 X373-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-INt 0 X373-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1403 X373-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-INt 0 X373-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-IN 0 z0=5 td=3.2ps
X373 X374-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-IN X373-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-INt X373-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-INt LSmitll_SPLITT

t1404 X374-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-INt 0 X374-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-IN 0 z0=5 td=3.7ps
t1405 X374-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-INt 0 X374-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-IN 0 z0=5 td=4.0ps
X374 X387-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-IN X374-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-INt X374-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-INt LSmitll_SPLITT

t1406 X375-LSmitll_SPLITT-OUT-X22-LSmitll_DFFT-INt 0 X375-LSmitll_SPLITT-OUT-X22-LSmitll_DFFT-IN 0 z0=5 td=3.3ps
t1407 X375-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-INt 0 X375-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
X375 X377-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-IN X375-LSmitll_SPLITT-OUT-X22-LSmitll_DFFT-INt X375-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-INt LSmitll_SPLITT

t1408 X376-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-INt 0 X376-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
t1409 X376-LSmitll_SPLITT-OUT-X187-LSmitll_AND2T-INt 0 X376-LSmitll_SPLITT-OUT-X187-LSmitll_AND2T-IN 0 z0=5 td=2.9ps
X376 X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-IN X376-LSmitll_SPLITT-OUT-X128-LSmitll_AND2T-INt X376-LSmitll_SPLITT-OUT-X187-LSmitll_AND2T-INt LSmitll_SPLITT

t1410 X377-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-INt 0 X377-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1411 X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-INt 0 X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X377 X380-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-IN X377-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-INt X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-INt LSmitll_SPLITT

t1412 X378-LSmitll_SPLITT-OUT-X129-LSmitll_DFFT-INt 0 X378-LSmitll_SPLITT-OUT-X129-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
t1413 X378-LSmitll_SPLITT-OUT-X131-LSmitll_DFFT-INt 0 X378-LSmitll_SPLITT-OUT-X131-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
X378 X379-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-IN X378-LSmitll_SPLITT-OUT-X129-LSmitll_DFFT-INt X378-LSmitll_SPLITT-OUT-X131-LSmitll_DFFT-INt LSmitll_SPLITT

t1414 X379-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-INt 0 X379-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
t1415 X379-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-INt 0 X379-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X379 X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-IN X379-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-INt X379-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-INt LSmitll_SPLITT

t1416 X380-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-INt 0 X380-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1417 X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-INt 0 X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
X380 X386-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-IN X380-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-INt X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-INt LSmitll_SPLITT

t1418 X381-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt 0 X381-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-IN 0 z0=5 td=4.7ps
t1419 X381-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-INt 0 X381-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-IN 0 z0=5 td=1.5ps
X381 X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-IN X381-LSmitll_SPLITT-OUT-X126-LSmitll_AND2T-INt X381-LSmitll_SPLITT-OUT-X158-LSmitll_AND2T-INt LSmitll_SPLITT

t1420 X382-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-INt 0 X382-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1421 X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-INt 0 X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X382 X385-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-IN X382-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-INt X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-INt LSmitll_SPLITT

t1422 X383-LSmitll_SPLITT-OUT-X127-LSmitll_DFFT-INt 0 X383-LSmitll_SPLITT-OUT-X127-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t1423 X383-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-INt 0 X383-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
X383 X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-IN X383-LSmitll_SPLITT-OUT-X127-LSmitll_DFFT-INt X383-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-INt LSmitll_SPLITT

t1424 X384-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-INt 0 X384-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1425 X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-INt 0 X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X384 X385-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-IN X384-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-INt X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-INt LSmitll_SPLITT

t1426 X385-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-INt 0 X385-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
t1427 X385-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-INt 0 X385-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X385 X386-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-IN X385-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-INt X385-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-INt LSmitll_SPLITT

t1428 X386-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-INt 0 X386-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-IN 0 z0=5 td=2.8ps
t1429 X386-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-INt 0 X386-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-IN 0 z0=5 td=4.5ps
X386 X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-IN X386-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-INt X386-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-INt LSmitll_SPLITT

t1430 X387-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-INt 0 X387-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t1431 X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-INt 0 X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-IN 0 z0=5 td=4.5ps
X387 X413-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-IN X387-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-INt X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-INt LSmitll_SPLITT

t1432 X388-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-INt 0 X388-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
t1433 X388-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-INt 0 X388-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-IN 0 z0=5 td=2.7ps
X388 X390-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-IN X388-LSmitll_SPLITT-OUT-X228-LSmitll_DFFT-INt X388-LSmitll_SPLITT-OUT-X239-LSmitll_AND2T-INt LSmitll_SPLITT

t1434 X389-LSmitll_SPLITT-OUT-X252-LSmitll_OR2T-INt 0 X389-LSmitll_SPLITT-OUT-X252-LSmitll_OR2T-IN 0 z0=5 td=1.1ps
t1435 X389-LSmitll_SPLITT-OUT-X253-LSmitll_DFFT-INt 0 X389-LSmitll_SPLITT-OUT-X253-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X389 X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-IN X389-LSmitll_SPLITT-OUT-X252-LSmitll_OR2T-INt X389-LSmitll_SPLITT-OUT-X253-LSmitll_DFFT-INt LSmitll_SPLITT

t1436 X390-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-INt 0 X390-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1437 X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-INt 0 X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X390 X393-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-IN X390-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-INt X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-INt LSmitll_SPLITT

t1438 X391-LSmitll_SPLITT-OUT-X184-LSmitll_AND2T-INt 0 X391-LSmitll_SPLITT-OUT-X184-LSmitll_AND2T-IN 0 z0=5 td=3.2ps
t1439 X391-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-INt 0 X391-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-IN 0 z0=5 td=1.3ps
X391 X392-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-IN X391-LSmitll_SPLITT-OUT-X184-LSmitll_AND2T-INt X391-LSmitll_SPLITT-OUT-X207-LSmitll_OR2T-INt LSmitll_SPLITT

t1440 X392-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-INt 0 X392-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1441 X392-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-INt 0 X392-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X392 X393-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-IN X392-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-INt X392-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-INt LSmitll_SPLITT

t1442 X393-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-INt 0 X393-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1443 X393-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-INt 0 X393-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X393 X399-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-IN X393-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-INt X393-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-INt LSmitll_SPLITT

t1444 X394-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt 0 X394-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1445 X394-LSmitll_SPLITT-OUT-X271-LSmitll_DFFT-INt 0 X394-LSmitll_SPLITT-OUT-X271-LSmitll_DFFT-IN 0 z0=5 td=4.7ps
X394 X395-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-IN X394-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt X394-LSmitll_SPLITT-OUT-X271-LSmitll_DFFT-INt LSmitll_SPLITT

t1446 X395-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-INt 0 X395-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1447 X395-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-INt 0 X395-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X395 X398-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-IN X395-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-INt X395-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-INt LSmitll_SPLITT

t1448 X396-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-INt 0 X396-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1449 X396-LSmitll_SPLITT-OUT-X205-LSmitll_DFFT-INt 0 X396-LSmitll_SPLITT-OUT-X205-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
X396 X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-IN X396-LSmitll_SPLITT-OUT-X191-LSmitll_AND2T-INt X396-LSmitll_SPLITT-OUT-X205-LSmitll_DFFT-INt LSmitll_SPLITT

t1450 X397-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-INt 0 X397-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
t1451 X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-INt 0 X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X397 X398-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-IN X397-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-INt X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-INt LSmitll_SPLITT

t1452 X398-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-INt 0 X398-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1453 X398-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-INt 0 X398-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-IN 0 z0=5 td=3.5ps
X398 X399-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-IN X398-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-INt X398-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-INt LSmitll_SPLITT

t1454 X399-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-INt 0 X399-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
t1455 X399-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-INt 0 X399-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X399 X412-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-IN X399-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-INt X399-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-INt LSmitll_SPLITT

t1456 X400-LSmitll_SPLITT-OUT-X141-LSmitll_XORT-INt 0 X400-LSmitll_SPLITT-OUT-X141-LSmitll_XORT-IN 0 z0=5 td=1.3ps
t1457 X400-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-INt 0 X400-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-IN 0 z0=5 td=1.9ps
X400 X402-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-IN X400-LSmitll_SPLITT-OUT-X141-LSmitll_XORT-INt X400-LSmitll_SPLITT-OUT-X156-LSmitll_AND2T-INt LSmitll_SPLITT

t1458 X401-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-INt 0 X401-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-IN 0 z0=5 td=0.9ps
t1459 X401-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-INt 0 X401-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
X401 X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-IN X401-LSmitll_SPLITT-OUT-X157-LSmitll_XORT-INt X401-LSmitll_SPLITT-OUT-X183-LSmitll_AND2T-INt LSmitll_SPLITT

t1460 X402-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-INt 0 X402-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
t1461 X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-INt 0 X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X402 X405-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-IN X402-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-INt X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-INt LSmitll_SPLITT

t1462 X403-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-INt 0 X403-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
t1463 X403-LSmitll_SPLITT-OUT-X125-LSmitll_DFFT-INt 0 X403-LSmitll_SPLITT-OUT-X125-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
X403 X404-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-IN X403-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-INt X403-LSmitll_SPLITT-OUT-X125-LSmitll_DFFT-INt LSmitll_SPLITT

t1464 X404-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-INt 0 X404-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
t1465 X404-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-INt 0 X404-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X404 X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-IN X404-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-INt X404-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-INt LSmitll_SPLITT

t1466 X405-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-INt 0 X405-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
t1467 X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-INt 0 X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
X405 X411-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-IN X405-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-INt X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-INt LSmitll_SPLITT

t1468 X406-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-INt 0 X406-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-IN 0 z0=5 td=5.1ps
t1469 X406-LSmitll_SPLITT-OUT-X200-LSmitll_OR2T-INt 0 X406-LSmitll_SPLITT-OUT-X200-LSmitll_OR2T-IN 0 z0=5 td=1.9ps
X406 X407-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-IN X406-LSmitll_SPLITT-OUT-X33-LSmitll_DFFT-INt X406-LSmitll_SPLITT-OUT-X200-LSmitll_OR2T-INt LSmitll_SPLITT

t1470 X407-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-INt 0 X407-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1471 X407-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-INt 0 X407-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X407 X410-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-IN X407-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-INt X407-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-INt LSmitll_SPLITT

t1472 X408-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-INt 0 X408-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
t1473 X408-LSmitll_SPLITT-OUT-X123-LSmitll_DFFT-INt 0 X408-LSmitll_SPLITT-OUT-X123-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
X408 X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-IN X408-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-INt X408-LSmitll_SPLITT-OUT-X123-LSmitll_DFFT-INt LSmitll_SPLITT

t1474 X409-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-INt 0 X409-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1475 X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-INt 0 X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X409 X410-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-IN X409-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-INt X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-INt LSmitll_SPLITT

t1476 X410-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-INt 0 X410-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
t1477 X410-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-INt 0 X410-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-IN 0 z0=5 td=3.5ps
X410 X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-IN X410-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-INt X410-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-INt LSmitll_SPLITT

t1478 X411-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-INt 0 X411-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1479 X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-INt 0 X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X411 X412-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-IN X411-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-INt X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-INt LSmitll_SPLITT

t1480 X412-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-INt 0 X412-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
t1481 X412-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-INt 0 X412-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-IN 0 z0=5 td=5.0ps
X412 X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-IN X412-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-INt X412-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-INt LSmitll_SPLITT

t1482 X413-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-INt 0 X413-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-IN 0 z0=5 td=4.7ps
t1483 X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-INt 0 X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-IN 0 z0=5 td=6.1ps
X413 X414-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-IN X413-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-INt X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-INt LSmitll_SPLITT

t1484 X414-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-INt 0 X414-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-IN 0 z0=5 td=5.2ps
t1485 X414-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-INt 0 X414-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-IN 0 z0=5 td=4.5ps
X414 X564-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-IN X414-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-INt X414-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-INt LSmitll_SPLITT

t1486 X415-LSmitll_SPLITT-OUT-X25-LSmitll_NOTT-INt 0 X415-LSmitll_SPLITT-OUT-X25-LSmitll_NOTT-IN 0 z0=5 td=1.6ps
t1487 X415-LSmitll_SPLITT-OUT-X76-LSmitll_OR2T-INt 0 X415-LSmitll_SPLITT-OUT-X76-LSmitll_OR2T-IN 0 z0=5 td=1.5ps
X415 X417-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-IN X415-LSmitll_SPLITT-OUT-X25-LSmitll_NOTT-INt X415-LSmitll_SPLITT-OUT-X76-LSmitll_OR2T-INt LSmitll_SPLITT

t1488 X416-LSmitll_SPLITT-OUT-X74-LSmitll_OR2T-INt 0 X416-LSmitll_SPLITT-OUT-X74-LSmitll_OR2T-IN 0 z0=5 td=1.0ps
t1489 X416-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-INt 0 X416-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-IN 0 z0=5 td=0.4ps
X416 X417-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-IN X416-LSmitll_SPLITT-OUT-X74-LSmitll_OR2T-INt X416-LSmitll_SPLITT-OUT-X77-LSmitll_DFFT-INt LSmitll_SPLITT

t1490 X417-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-INt 0 X417-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
t1491 X417-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-INt 0 X417-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X417 X420-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-IN X417-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-INt X417-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-INt LSmitll_SPLITT

t1492 X418-LSmitll_SPLITT-OUT-X115-LSmitll_NDROT-INt 0 X418-LSmitll_SPLITT-OUT-X115-LSmitll_NDROT-IN 0 z0=5 td=1.9ps
t1493 X418-LSmitll_SPLITT-OUT-X116-LSmitll_AND2T-INt 0 X418-LSmitll_SPLITT-OUT-X116-LSmitll_AND2T-IN 0 z0=5 td=1.3ps
X418 X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-IN X418-LSmitll_SPLITT-OUT-X115-LSmitll_NDROT-INt X418-LSmitll_SPLITT-OUT-X116-LSmitll_AND2T-INt LSmitll_SPLITT

t1494 X419-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-INt 0 X419-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1495 X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-INt 0 X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X419 X420-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-IN X419-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-INt X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-INt LSmitll_SPLITT

t1496 X420-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-INt 0 X420-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1497 X420-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-INt 0 X420-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X420 X427-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-IN X420-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-INt X420-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-INt LSmitll_SPLITT

t1498 X421-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-INt 0 X421-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-IN 0 z0=5 td=0.4ps
t1499 X421-LSmitll_SPLITT-OUT-X59-LSmitll_AND2T-INt 0 X421-LSmitll_SPLITT-OUT-X59-LSmitll_AND2T-IN 0 z0=5 td=1.4ps
X421 X423-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-IN X421-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-INt X421-LSmitll_SPLITT-OUT-X59-LSmitll_AND2T-INt LSmitll_SPLITT

t1500 X422-LSmitll_SPLITT-OUT-X2-LSmitll_DFFT-INt 0 X422-LSmitll_SPLITT-OUT-X2-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
t1501 X422-LSmitll_SPLITT-OUT-X60-LSmitll_AND2T-INt 0 X422-LSmitll_SPLITT-OUT-X60-LSmitll_AND2T-IN 0 z0=5 td=0.4ps
X422 X423-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-IN X422-LSmitll_SPLITT-OUT-X2-LSmitll_DFFT-INt X422-LSmitll_SPLITT-OUT-X60-LSmitll_AND2T-INt LSmitll_SPLITT

t1502 X423-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-INt 0 X423-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
t1503 X423-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-INt 0 X423-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X423 X426-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-IN X423-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-INt X423-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-INt LSmitll_SPLITT

t1504 X424-LSmitll_SPLITT-OUT-X91-LSmitll_NDROT-INt 0 X424-LSmitll_SPLITT-OUT-X91-LSmitll_NDROT-IN 0 z0=5 td=3.8ps
t1505 X424-LSmitll_SPLITT-OUT-X309-LSmitll_DFFT-INt 0 X424-LSmitll_SPLITT-OUT-X309-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X424 X425-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-IN X424-LSmitll_SPLITT-OUT-X91-LSmitll_NDROT-INt X424-LSmitll_SPLITT-OUT-X309-LSmitll_DFFT-INt LSmitll_SPLITT

t1506 X425-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-INt 0 X425-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
t1507 X425-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-INt 0 X425-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X425 X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-IN X425-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-INt X425-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-INt LSmitll_SPLITT

t1508 X426-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-INt 0 X426-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1509 X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-INt 0 X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X426 X427-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-IN X426-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-INt X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-INt LSmitll_SPLITT

t1510 X427-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-INt 0 X427-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1511 X427-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-INt 0 X427-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X427 X440-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-IN X427-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-INt X427-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-INt LSmitll_SPLITT

t1512 X428-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-INt 0 X428-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t1513 X428-LSmitll_SPLITT-OUT-X280-LSmitll_OR2T-INt 0 X428-LSmitll_SPLITT-OUT-X280-LSmitll_OR2T-IN 0 z0=5 td=0.7ps
X428 X430-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-IN X428-LSmitll_SPLITT-OUT-X86-LSmitll_AND2T-INt X428-LSmitll_SPLITT-OUT-X280-LSmitll_OR2T-INt LSmitll_SPLITT

t1514 X429-LSmitll_SPLITT-OUT-X85-LSmitll_NDROT-INt 0 X429-LSmitll_SPLITT-OUT-X85-LSmitll_NDROT-IN 0 z0=5 td=0.6ps
t1515 X429-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-INt 0 X429-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
X429 X430-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-IN X429-LSmitll_SPLITT-OUT-X85-LSmitll_NDROT-INt X429-LSmitll_SPLITT-OUT-X92-LSmitll_AND2T-INt LSmitll_SPLITT

t1516 X430-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-INt 0 X430-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-IN 0 z0=5 td=2.8ps
t1517 X430-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-INt 0 X430-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X430 X433-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-IN X430-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-INt X430-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-INt LSmitll_SPLITT

t1518 X431-LSmitll_SPLITT-OUT-X282-LSmitll_OR2T-INt 0 X431-LSmitll_SPLITT-OUT-X282-LSmitll_OR2T-IN 0 z0=5 td=2.8ps
t1519 X431-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-INt 0 X431-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
X431 X432-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-IN X431-LSmitll_SPLITT-OUT-X282-LSmitll_OR2T-INt X431-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-INt LSmitll_SPLITT

t1520 X432-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-INt 0 X432-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1521 X432-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-INt 0 X432-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X432 X433-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-IN X432-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-INt X432-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-INt LSmitll_SPLITT

t1522 X433-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-INt 0 X433-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1523 X433-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-INt 0 X433-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X433 X439-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-IN X433-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-INt X433-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-INt LSmitll_SPLITT

t1524 X434-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-INt 0 X434-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-IN 0 z0=5 td=0.4ps
t1525 X434-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-INt 0 X434-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
X434 X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-IN X434-LSmitll_SPLITT-OUT-X89-LSmitll_AND2T-INt X434-LSmitll_SPLITT-OUT-X276-LSmitll_DFFT-INt LSmitll_SPLITT

t1526 X435-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-INt 0 X435-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1527 X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-INt 0 X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X435 X438-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-IN X435-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-INt X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-INt LSmitll_SPLITT

t1528 X436-LSmitll_SPLITT-OUT-X88-LSmitll_NDROT-INt 0 X436-LSmitll_SPLITT-OUT-X88-LSmitll_NDROT-IN 0 z0=5 td=0.9ps
t1529 X436-LSmitll_SPLITT-OUT-X233-LSmitll_DFFT-INt 0 X436-LSmitll_SPLITT-OUT-X233-LSmitll_DFFT-IN 0 z0=5 td=5.6ps
X436 X437-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-IN X436-LSmitll_SPLITT-OUT-X88-LSmitll_NDROT-INt X436-LSmitll_SPLITT-OUT-X233-LSmitll_DFFT-INt LSmitll_SPLITT

t1530 X437-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-INt 0 X437-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1531 X437-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-INt 0 X437-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X437 X438-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-IN X437-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-INt X437-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-INt LSmitll_SPLITT

t1532 X438-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-INt 0 X438-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
t1533 X438-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-INt 0 X438-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X438 X439-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-IN X438-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-INt X438-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-INt LSmitll_SPLITT

t1534 X439-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-INt 0 X439-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
t1535 X439-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-INt 0 X439-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X439 X440-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-IN X439-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-INt X439-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-INt LSmitll_SPLITT

t1536 X440-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-INt 0 X440-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-IN 0 z0=5 td=5.8ps
t1537 X440-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-INt 0 X440-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X440 X466-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-IN X440-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-INt X440-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-INt LSmitll_SPLITT

t1538 X441-LSmitll_SPLITT-OUT-X23-LSmitll_NOTT-INt 0 X441-LSmitll_SPLITT-OUT-X23-LSmitll_NOTT-IN 0 z0=5 td=1.8ps
t1539 X441-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-INt 0 X441-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X441 X443-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-IN X441-LSmitll_SPLITT-OUT-X23-LSmitll_NOTT-INt X441-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-INt LSmitll_SPLITT

t1540 X442-LSmitll_SPLITT-OUT-X57-LSmitll_AND2T-INt 0 X442-LSmitll_SPLITT-OUT-X57-LSmitll_AND2T-IN 0 z0=5 td=1.4ps
t1541 X442-LSmitll_SPLITT-OUT-X58-LSmitll_AND2T-INt 0 X442-LSmitll_SPLITT-OUT-X58-LSmitll_AND2T-IN 0 z0=5 td=0.5ps
X442 X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-IN X442-LSmitll_SPLITT-OUT-X57-LSmitll_AND2T-INt X442-LSmitll_SPLITT-OUT-X58-LSmitll_AND2T-INt LSmitll_SPLITT

t1542 X443-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-INt 0 X443-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1543 X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-INt 0 X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X443 X446-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-IN X443-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-INt X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-INt LSmitll_SPLITT

t1544 X444-LSmitll_SPLITT-OUT-X39-LSmitll_DFFT-INt 0 X444-LSmitll_SPLITT-OUT-X39-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
t1545 X444-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-INt 0 X444-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
X444 X445-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-IN X444-LSmitll_SPLITT-OUT-X39-LSmitll_DFFT-INt X444-LSmitll_SPLITT-OUT-X78-LSmitll_DFFT-INt LSmitll_SPLITT

t1546 X445-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-INt 0 X445-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1547 X445-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-INt 0 X445-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X445 X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-IN X445-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-INt X445-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-INt LSmitll_SPLITT

t1548 X446-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-INt 0 X446-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1549 X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-INt 0 X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
X446 X452-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-IN X446-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-INt X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-INt LSmitll_SPLITT

t1550 X447-LSmitll_SPLITT-OUT-X73-LSmitll_OR2T-INt 0 X447-LSmitll_SPLITT-OUT-X73-LSmitll_OR2T-IN 0 z0=5 td=2.1ps
t1551 X447-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-INt 0 X447-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
X447 X448-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-IN X447-LSmitll_SPLITT-OUT-X73-LSmitll_OR2T-INt X447-LSmitll_SPLITT-OUT-X303-LSmitll_DFFT-INt LSmitll_SPLITT

t1552 X448-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-INt 0 X448-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
t1553 X448-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-INt 0 X448-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
X448 X451-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-IN X448-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-INt X448-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-INt LSmitll_SPLITT

t1554 X449-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-INt 0 X449-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1555 X449-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-INt 0 X449-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X449 X450-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-IN X449-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-INt X449-LSmitll_SPLITT-OUT-X298-LSmitll_DFFT-INt LSmitll_SPLITT

t1556 X450-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-INt 0 X450-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1557 X450-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-INt 0 X450-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X450 X451-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-IN X450-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-INt X450-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-INt LSmitll_SPLITT

t1558 X451-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-INt 0 X451-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1559 X451-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-INt 0 X451-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X451 X452-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-IN X451-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-INt X451-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-INt LSmitll_SPLITT

t1560 X452-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-INt 0 X452-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
t1561 X452-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-INt 0 X452-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X452 X465-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-IN X452-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-INt X452-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-INt LSmitll_SPLITT

t1562 X453-LSmitll_SPLITT-OUT-X267-LSmitll_DFFT-INt 0 X453-LSmitll_SPLITT-OUT-X267-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
t1563 X453-LSmitll_SPLITT-OUT-X288-LSmitll_XORT-INt 0 X453-LSmitll_SPLITT-OUT-X288-LSmitll_XORT-IN 0 z0=5 td=2.0ps
X453 X455-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-IN X453-LSmitll_SPLITT-OUT-X267-LSmitll_DFFT-INt X453-LSmitll_SPLITT-OUT-X288-LSmitll_XORT-INt LSmitll_SPLITT

t1564 X454-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-INt 0 X454-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-IN 0 z0=5 td=1.3ps
t1565 X454-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-INt 0 X454-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
X454 X455-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-IN X454-LSmitll_SPLITT-OUT-X95-LSmitll_AND2T-INt X454-LSmitll_SPLITT-OUT-X277-LSmitll_DFFT-INt LSmitll_SPLITT

t1566 X455-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-INt 0 X455-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1567 X455-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-INt 0 X455-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X455 X458-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-IN X455-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-INt X455-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-INt LSmitll_SPLITT

t1568 X456-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-INt 0 X456-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
t1569 X456-LSmitll_SPLITT-OUT-X270-LSmitll_DFFT-INt 0 X456-LSmitll_SPLITT-OUT-X270-LSmitll_DFFT-IN 0 z0=5 td=2.7ps
X456 X457-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-IN X456-LSmitll_SPLITT-OUT-X261-LSmitll_DFFT-INt X456-LSmitll_SPLITT-OUT-X270-LSmitll_DFFT-INt LSmitll_SPLITT

t1570 X457-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-INt 0 X457-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1571 X457-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-INt 0 X457-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X457 X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-IN X457-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-INt X457-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-INt LSmitll_SPLITT

t1572 X458-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-INt 0 X458-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1573 X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-INt 0 X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X458 X464-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-IN X458-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-INt X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-INt LSmitll_SPLITT

t1574 X459-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-INt 0 X459-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-IN 0 z0=5 td=1.8ps
t1575 X459-LSmitll_SPLITT-OUT-X283-LSmitll_DFFT-INt 0 X459-LSmitll_SPLITT-OUT-X283-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
X459 X460-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-IN X459-LSmitll_SPLITT-OUT-X262-LSmitll_DFFT-INt X459-LSmitll_SPLITT-OUT-X283-LSmitll_DFFT-INt LSmitll_SPLITT

t1576 X460-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-INt 0 X460-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-IN 0 z0=5 td=2.8ps
t1577 X460-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-INt 0 X460-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X460 X463-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-IN X460-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-INt X460-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-INt LSmitll_SPLITT

t1578 X461-LSmitll_SPLITT-OUT-X291-LSmitll_XORT-INt 0 X461-LSmitll_SPLITT-OUT-X291-LSmitll_XORT-IN 0 z0=5 td=1.7ps
t1579 X461-LSmitll_SPLITT-OUT-X296-LSmitll_XORT-INt 0 X461-LSmitll_SPLITT-OUT-X296-LSmitll_XORT-IN 0 z0=5 td=1.7ps
X461 X462-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-IN X461-LSmitll_SPLITT-OUT-X291-LSmitll_XORT-INt X461-LSmitll_SPLITT-OUT-X296-LSmitll_XORT-INt LSmitll_SPLITT

t1580 X462-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-INt 0 X462-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1581 X462-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-INt 0 X462-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X462 X463-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-IN X462-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-INt X462-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-INt LSmitll_SPLITT

t1582 X463-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-INt 0 X463-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1583 X463-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-INt 0 X463-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X463 X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-IN X463-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-INt X463-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-INt LSmitll_SPLITT

t1584 X464-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-INt 0 X464-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1585 X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-INt 0 X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X464 X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-IN X464-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-INt X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-INt LSmitll_SPLITT

t1586 X465-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-INt 0 X465-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1587 X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-INt 0 X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
X465 X466-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-IN X465-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-INt X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-INt LSmitll_SPLITT

t1588 X466-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-INt 0 X466-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-IN 0 z0=5 td=4.6ps
t1589 X466-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-INt 0 X466-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-IN 0 z0=5 td=4.0ps
X466 X518-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-IN X466-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-INt X466-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-INt LSmitll_SPLITT

t1590 X467-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-INt 0 X467-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
t1591 X467-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-INt 0 X467-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
X467 X469-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-IN X467-LSmitll_SPLITT-OUT-X231-LSmitll_AND2T-INt X467-LSmitll_SPLITT-OUT-X274-LSmitll_DFFT-INt LSmitll_SPLITT

t1592 X468-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-INt 0 X468-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t1593 X468-LSmitll_SPLITT-OUT-X268-LSmitll_DFFT-INt 0 X468-LSmitll_SPLITT-OUT-X268-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
X468 X469-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-IN X468-LSmitll_SPLITT-OUT-X235-LSmitll_AND2T-INt X468-LSmitll_SPLITT-OUT-X268-LSmitll_DFFT-INt LSmitll_SPLITT

t1594 X469-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-INt 0 X469-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t1595 X469-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-INt 0 X469-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X469 X472-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-IN X469-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-INt X469-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-INt LSmitll_SPLITT

t1596 X470-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-INt 0 X470-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-IN 0 z0=5 td=0.8ps
t1597 X470-LSmitll_SPLITT-OUT-X203-LSmitll_DFFT-INt 0 X470-LSmitll_SPLITT-OUT-X203-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
X470 X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-IN X470-LSmitll_SPLITT-OUT-X188-LSmitll_AND2T-INt X470-LSmitll_SPLITT-OUT-X203-LSmitll_DFFT-INt LSmitll_SPLITT

t1598 X471-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-INt 0 X471-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
t1599 X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-INt 0 X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X471 X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-IN X471-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-INt X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-INt LSmitll_SPLITT

t1600 X472-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-INt 0 X472-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
t1601 X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-INt 0 X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
X472 X478-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-IN X472-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-INt X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-INt LSmitll_SPLITT

t1602 X473-LSmitll_SPLITT-OUT-X248-LSmitll_DFFT-INt 0 X473-LSmitll_SPLITT-OUT-X248-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
t1603 X473-LSmitll_SPLITT-OUT-X250-LSmitll_DFFT-INt 0 X473-LSmitll_SPLITT-OUT-X250-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X473 X474-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-IN X473-LSmitll_SPLITT-OUT-X248-LSmitll_DFFT-INt X473-LSmitll_SPLITT-OUT-X250-LSmitll_DFFT-INt LSmitll_SPLITT

t1604 X474-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-INt 0 X474-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1605 X474-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-INt 0 X474-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X474 X477-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-IN X474-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-INt X474-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-INt LSmitll_SPLITT

t1606 X475-LSmitll_SPLITT-OUT-X112-LSmitll_NDROT-INt 0 X475-LSmitll_SPLITT-OUT-X112-LSmitll_NDROT-IN 0 z0=5 td=1.1ps
t1607 X475-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-INt 0 X475-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X475 X476-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-IN X475-LSmitll_SPLITT-OUT-X112-LSmitll_NDROT-INt X475-LSmitll_SPLITT-OUT-X204-LSmitll_OR2T-INt LSmitll_SPLITT

t1608 X476-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-INt 0 X476-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1609 X476-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-INt 0 X476-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X476 X477-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-IN X476-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-INt X476-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-INt LSmitll_SPLITT

t1610 X477-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-INt 0 X477-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1611 X477-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-INt 0 X477-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X477 X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-IN X477-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-INt X477-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-INt LSmitll_SPLITT

t1612 X478-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-INt 0 X478-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
t1613 X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-INt 0 X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X478 X491-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-IN X478-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-INt X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-INt LSmitll_SPLITT

t1614 X479-LSmitll_SPLITT-OUT-X145-LSmitll_XORT-INt 0 X479-LSmitll_SPLITT-OUT-X145-LSmitll_XORT-IN 0 z0=5 td=2.0ps
t1615 X479-LSmitll_SPLITT-OUT-X193-LSmitll_AND2T-INt 0 X479-LSmitll_SPLITT-OUT-X193-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X479 X481-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-IN X479-LSmitll_SPLITT-OUT-X145-LSmitll_XORT-INt X479-LSmitll_SPLITT-OUT-X193-LSmitll_AND2T-INt LSmitll_SPLITT

t1616 X480-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt 0 X480-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-IN 0 z0=5 td=4.3ps
t1617 X480-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-INt 0 X480-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-IN 0 z0=5 td=2.4ps
X480 X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-IN X480-LSmitll_SPLITT-OUT-X132-LSmitll_AND2T-INt X480-LSmitll_SPLITT-OUT-X208-LSmitll_OR2T-INt LSmitll_SPLITT

t1618 X481-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-INt 0 X481-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1619 X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-INt 0 X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X481 X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-IN X481-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-INt X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-INt LSmitll_SPLITT

t1620 X482-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-INt 0 X482-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-IN 0 z0=5 td=4.3ps
t1621 X482-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-INt 0 X482-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-IN 0 z0=5 td=0.4ps
X482 X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-IN X482-LSmitll_SPLITT-OUT-X118-LSmitll_AND2T-INt X482-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-INt LSmitll_SPLITT

t1622 X483-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-INt 0 X483-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1623 X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-INt 0 X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X483 X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-IN X483-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-INt X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-INt LSmitll_SPLITT

t1624 X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-INt 0 X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-IN 0 z0=5 td=0.5ps
t1625 X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-INt 0 X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-IN 0 z0=5 td=3.4ps
X484 X490-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-IN X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-INt X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-INt LSmitll_SPLITT

t1626 X485-LSmitll_SPLITT-OUT-X147-LSmitll_XORT-INt 0 X485-LSmitll_SPLITT-OUT-X147-LSmitll_XORT-IN 0 z0=5 td=2.7ps
t1627 X485-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-INt 0 X485-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
X485 X486-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-IN X485-LSmitll_SPLITT-OUT-X147-LSmitll_XORT-INt X485-LSmitll_SPLITT-OUT-X192-LSmitll_AND2T-INt LSmitll_SPLITT

t1628 X486-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-INt 0 X486-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1629 X486-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-INt 0 X486-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X486 X489-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-IN X486-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-INt X486-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-INt LSmitll_SPLITT

t1630 X487-LSmitll_SPLITT-OUT-X68-LSmitll_DFFT-INt 0 X487-LSmitll_SPLITT-OUT-X68-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
t1631 X487-LSmitll_SPLITT-OUT-X119-LSmitll_DFFT-INt 0 X487-LSmitll_SPLITT-OUT-X119-LSmitll_DFFT-IN 0 z0=5 td=3.3ps
X487 X488-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-IN X487-LSmitll_SPLITT-OUT-X68-LSmitll_DFFT-INt X487-LSmitll_SPLITT-OUT-X119-LSmitll_DFFT-INt LSmitll_SPLITT

t1632 X488-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-INt 0 X488-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
t1633 X488-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-INt 0 X488-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X488 X489-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-IN X488-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-INt X488-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-INt LSmitll_SPLITT

t1634 X489-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-INt 0 X489-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-IN 0 z0=5 td=6.1ps
t1635 X489-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-INt 0 X489-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X489 X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-IN X489-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-INt X489-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-INt LSmitll_SPLITT

t1636 X490-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-INt 0 X490-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
t1637 X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-INt 0 X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X490 X491-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-IN X490-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-INt X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-INt LSmitll_SPLITT

t1638 X491-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-INt 0 X491-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
t1639 X491-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-INt 0 X491-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X491 X517-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-IN X491-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-INt X491-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-INt LSmitll_SPLITT

t1640 X492-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt 0 X492-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
t1641 X492-LSmitll_SPLITT-OUT-X294-LSmitll_DFFT-INt 0 X492-LSmitll_SPLITT-OUT-X294-LSmitll_DFFT-IN 0 z0=5 td=7.2ps
X492 X494-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-IN X492-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt X492-LSmitll_SPLITT-OUT-X294-LSmitll_DFFT-INt LSmitll_SPLITT

t1642 X493-LSmitll_SPLITT-OUT-X232-LSmitll_DFFT-INt 0 X493-LSmitll_SPLITT-OUT-X232-LSmitll_DFFT-IN 0 z0=5 td=2.0ps
t1643 X493-LSmitll_SPLITT-OUT-X249-LSmitll_OR2T-INt 0 X493-LSmitll_SPLITT-OUT-X249-LSmitll_OR2T-IN 0 z0=5 td=2.4ps
X493 X494-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-IN X493-LSmitll_SPLITT-OUT-X232-LSmitll_DFFT-INt X493-LSmitll_SPLITT-OUT-X249-LSmitll_OR2T-INt LSmitll_SPLITT

t1644 X494-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-INt 0 X494-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1645 X494-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-INt 0 X494-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X494 X497-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-IN X494-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-INt X494-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-INt LSmitll_SPLITT

t1646 X495-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-INt 0 X495-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1647 X495-LSmitll_SPLITT-OUT-X308-LSmitll_DFFT-INt 0 X495-LSmitll_SPLITT-OUT-X308-LSmitll_DFFT-IN 0 z0=5 td=3.4ps
X495 X496-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-IN X495-LSmitll_SPLITT-OUT-X189-LSmitll_AND2T-INt X495-LSmitll_SPLITT-OUT-X308-LSmitll_DFFT-INt LSmitll_SPLITT

t1648 X496-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-INt 0 X496-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t1649 X496-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-INt 0 X496-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X496 X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-IN X496-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-INt X496-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-INt LSmitll_SPLITT

t1650 X497-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-INt 0 X497-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1651 X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-INt 0 X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X497 X503-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-IN X497-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-INt X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-INt LSmitll_SPLITT

t1652 X498-LSmitll_SPLITT-OUT-X110-LSmitll_AND2T-INt 0 X498-LSmitll_SPLITT-OUT-X110-LSmitll_AND2T-IN 0 z0=5 td=0.7ps
t1653 X498-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-INt 0 X498-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-IN 0 z0=5 td=5.2ps
X498 X499-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-IN X498-LSmitll_SPLITT-OUT-X110-LSmitll_AND2T-INt X498-LSmitll_SPLITT-OUT-X237-LSmitll_DFFT-INt LSmitll_SPLITT

t1654 X499-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-INt 0 X499-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1655 X499-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-INt 0 X499-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X499 X502-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-IN X499-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-INt X499-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-INt LSmitll_SPLITT

t1656 X500-LSmitll_SPLITT-OUT-X109-LSmitll_NDROT-INt 0 X500-LSmitll_SPLITT-OUT-X109-LSmitll_NDROT-IN 0 z0=5 td=2.4ps
t1657 X500-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-INt 0 X500-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-IN 0 z0=5 td=3.3ps
X500 X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-IN X500-LSmitll_SPLITT-OUT-X109-LSmitll_NDROT-INt X500-LSmitll_SPLITT-OUT-X160-LSmitll_AND2T-INt LSmitll_SPLITT

t1658 X501-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-INt 0 X501-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1659 X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-INt 0 X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X501 X502-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-IN X501-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-INt X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-INt LSmitll_SPLITT

t1660 X502-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-INt 0 X502-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-IN 0 z0=5 td=4.2ps
t1661 X502-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-INt 0 X502-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
X502 X503-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-IN X502-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-INt X502-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-INt LSmitll_SPLITT

t1662 X503-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-INt 0 X503-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1663 X503-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-INt 0 X503-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-IN 0 z0=5 td=4.1ps
X503 X516-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-IN X503-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-INt X503-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-INt LSmitll_SPLITT

t1664 X504-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt 0 X504-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-IN 0 z0=5 td=0.5ps
t1665 X504-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-INt 0 X504-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
X504 X506-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-IN X504-LSmitll_SPLITT-OUT-X122-LSmitll_AND2T-INt X504-LSmitll_SPLITT-OUT-X162-LSmitll_AND2T-INt LSmitll_SPLITT

t1666 X505-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-INt 0 X505-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-IN 0 z0=5 td=3.5ps
t1667 X505-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-INt 0 X505-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-IN 0 z0=5 td=1.7ps
X505 X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-IN X505-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-INt X505-LSmitll_SPLITT-OUT-X163-LSmitll_XORT-INt LSmitll_SPLITT

t1668 X506-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-INt 0 X506-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1669 X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-INt 0 X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X506 X509-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-IN X506-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-INt X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-INt LSmitll_SPLITT

t1670 X507-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-INt 0 X507-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-IN 0 z0=5 td=1.4ps
t1671 X507-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-INt 0 X507-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
X507 X508-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-IN X507-LSmitll_SPLITT-OUT-X66-LSmitll_DFFT-INt X507-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-INt LSmitll_SPLITT

t1672 X508-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-INt 0 X508-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1673 X508-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-INt 0 X508-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X508 X509-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-IN X508-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-INt X508-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-INt LSmitll_SPLITT

t1674 X509-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-INt 0 X509-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1675 X509-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-INt 0 X509-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X509 X515-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-IN X509-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-INt X509-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-INt LSmitll_SPLITT

t1676 X510-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt 0 X510-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-IN 0 z0=5 td=3.1ps
t1677 X510-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-INt 0 X510-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-IN 0 z0=5 td=2.8ps
X510 X511-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-IN X510-LSmitll_SPLITT-OUT-X124-LSmitll_AND2T-INt X510-LSmitll_SPLITT-OUT-X161-LSmitll_XORT-INt LSmitll_SPLITT

t1678 X511-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-INt 0 X511-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1679 X511-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-INt 0 X511-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X511 X514-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-IN X511-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-INt X511-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-INt LSmitll_SPLITT

t1680 X512-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-INt 0 X512-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
t1681 X512-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-INt 0 X512-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X512 X513-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-IN X512-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-INt X512-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-INt LSmitll_SPLITT

t1682 X513-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-INt 0 X513-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1683 X513-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-INt 0 X513-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X513 X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-IN X513-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-INt X513-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-INt LSmitll_SPLITT

t1684 X514-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-INt 0 X514-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
t1685 X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-INt 0 X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
X514 X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-IN X514-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-INt X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-INt LSmitll_SPLITT

t1686 X515-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-INt 0 X515-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1687 X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-INt 0 X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X515 X516-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-IN X515-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-INt X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-INt LSmitll_SPLITT

t1688 X516-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-INt 0 X516-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
t1689 X516-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-INt 0 X516-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-IN 0 z0=5 td=3.7ps
X516 X517-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-IN X516-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-INt X516-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-INt LSmitll_SPLITT

t1690 X517-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-INt 0 X517-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
t1691 X517-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-INt 0 X517-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
X517 X518-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-IN X517-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-INt X517-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-INt LSmitll_SPLITT

t1692 X518-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-INt 0 X518-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-IN 0 z0=5 td=8.0ps
t1693 X518-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-INt 0 X518-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-IN 0 z0=5 td=7.2ps
X518 X564-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-IN X518-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-INt X518-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-INt LSmitll_SPLITT

t1694 X519-LSmitll_SPLITT-OUT-X1-LSmitll_DFFT-INt 0 X519-LSmitll_SPLITT-OUT-X1-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1695 X519-SPLITT-OUT-R-INt 0 X519-SPLITT-OUT-R-IN 0 z0=5 td=9.9ps
X519 X448-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-IN X519-LSmitll_SPLITT-OUT-X1-LSmitll_DFFT-INt X519-SPLITT-OUT-R-INt LSmitll_SPLITT

t1696 X520-LSmitll_SPLITT-OUT-X7-LSmitll_DFFT-INt 0 X520-LSmitll_SPLITT-OUT-X7-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1697 X520-SPLITT-OUT-R-INt 0 X520-SPLITT-OUT-R-IN 0 z0=5 td=10.2ps
X520 X343-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-IN X520-LSmitll_SPLITT-OUT-X7-LSmitll_DFFT-INt X520-SPLITT-OUT-R-INt LSmitll_SPLITT

t1698 X521-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-INt 0 X521-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1699 X521-SPLITT-OUT-R-INt 0 X521-SPLITT-OUT-R-IN 0 z0=5 td=10.0ps
X521 X513-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-IN X521-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-INt X521-SPLITT-OUT-R-INt LSmitll_SPLITT

t1700 X522-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-INt 0 X522-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1701 X522-SPLITT-OUT-R-INt 0 X522-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X522 X483-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-IN X522-LSmitll_SPLITT-OUT-X34-LSmitll_DFFT-INt X522-SPLITT-OUT-R-INt LSmitll_SPLITT

t1702 X523-LSmitll_SPLITT-OUT-X63-LSmitll_AND2T-INt 0 X523-LSmitll_SPLITT-OUT-X63-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
t1703 X523-SPLITT-OUT-R-INt 0 X523-SPLITT-OUT-R-IN 0 z0=5 td=9.7ps
X523 X345-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-IN X523-LSmitll_SPLITT-OUT-X63-LSmitll_AND2T-INt X523-SPLITT-OUT-R-INt LSmitll_SPLITT

t1704 X524-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-INt 0 X524-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1705 X524-SPLITT-OUT-R-INt 0 X524-SPLITT-OUT-R-IN 0 z0=5 td=10.2ps
X524 X384-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-IN X524-LSmitll_SPLITT-OUT-X65-LSmitll_DFFT-INt X524-SPLITT-OUT-R-INt LSmitll_SPLITT

t1706 X525-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-INt 0 X525-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1707 X525-SPLITT-OUT-R-INt 0 X525-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X525 X404-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-IN X525-LSmitll_SPLITT-OUT-X67-LSmitll_DFFT-INt X525-SPLITT-OUT-R-INt LSmitll_SPLITT

t1708 X526-LSmitll_SPLITT-OUT-X80-LSmitll_DFFT-INt 0 X526-LSmitll_SPLITT-OUT-X80-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1709 X526-SPLITT-OUT-R-INt 0 X526-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X526 X314-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-IN X526-LSmitll_SPLITT-OUT-X80-LSmitll_DFFT-INt X526-SPLITT-OUT-R-INt LSmitll_SPLITT

t1710 X527-LSmitll_SPLITT-OUT-X94-LSmitll_NDROT-INt 0 X527-LSmitll_SPLITT-OUT-X94-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
t1711 X527-SPLITT-OUT-R-INt 0 X527-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X527 X450-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-IN X527-LSmitll_SPLITT-OUT-X94-LSmitll_NDROT-INt X527-SPLITT-OUT-R-INt LSmitll_SPLITT

t1712 X528-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-INt 0 X528-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
t1713 X528-SPLITT-OUT-R-INt 0 X528-SPLITT-OUT-R-IN 0 z0=5 td=10.0ps
X528 X330-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-IN X528-LSmitll_SPLITT-OUT-X98-LSmitll_AND2T-INt X528-SPLITT-OUT-R-INt LSmitll_SPLITT

t1714 X529-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt 0 X529-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
t1715 X529-SPLITT-OUT-R-INt 0 X529-SPLITT-OUT-R-IN 0 z0=5 td=9.9ps
X529 X320-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-IN X529-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt X529-SPLITT-OUT-R-INt LSmitll_SPLITT

t1716 X530-LSmitll_SPLITT-OUT-X106-LSmitll_NDROT-INt 0 X530-LSmitll_SPLITT-OUT-X106-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
t1717 X530-SPLITT-OUT-R-INt 0 X530-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X530 X340-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-IN X530-LSmitll_SPLITT-OUT-X106-LSmitll_NDROT-INt X530-SPLITT-OUT-R-INt LSmitll_SPLITT

t1718 X531-LSmitll_SPLITT-OUT-X113-LSmitll_AND2T-INt 0 X531-LSmitll_SPLITT-OUT-X113-LSmitll_AND2T-IN 0 z0=5 td=0.8ps
t1719 X531-SPLITT-OUT-R-INt 0 X531-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X531 X476-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-IN X531-LSmitll_SPLITT-OUT-X113-LSmitll_AND2T-INt X531-SPLITT-OUT-R-INt LSmitll_SPLITT

t1720 X532-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt 0 X532-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
t1721 X532-SPLITT-OUT-R-INt 0 X532-SPLITT-OUT-R-IN 0 z0=5 td=9.5ps
X532 X409-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-IN X532-LSmitll_SPLITT-OUT-X120-LSmitll_AND2T-INt X532-SPLITT-OUT-R-INt LSmitll_SPLITT

t1722 X533-LSmitll_SPLITT-OUT-X121-LSmitll_DFFT-INt 0 X533-LSmitll_SPLITT-OUT-X121-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1723 X533-SPLITT-OUT-R-INt 0 X533-SPLITT-OUT-R-IN 0 z0=5 td=10.5ps
X533 X488-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-IN X533-LSmitll_SPLITT-OUT-X121-LSmitll_DFFT-INt X533-SPLITT-OUT-R-INt LSmitll_SPLITT

t1724 X534-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt 0 X534-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-IN 0 z0=5 td=0.8ps
t1725 X534-SPLITT-OUT-R-INt 0 X534-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X534 X407-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-IN X534-LSmitll_SPLITT-OUT-X130-LSmitll_AND2T-INt X534-SPLITT-OUT-R-INt LSmitll_SPLITT

t1726 X535-LSmitll_SPLITT-OUT-X133-LSmitll_DFFT-INt 0 X535-LSmitll_SPLITT-OUT-X133-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1727 X535-SPLITT-OUT-R-INt 0 X535-SPLITT-OUT-R-IN 0 z0=5 td=9.5ps
X535 X511-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-IN X535-LSmitll_SPLITT-OUT-X133-LSmitll_DFFT-INt X535-SPLITT-OUT-R-INt LSmitll_SPLITT

t1728 X536-LSmitll_SPLITT-OUT-X134-LSmitll_DFFT-INt 0 X536-LSmitll_SPLITT-OUT-X134-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1729 X536-SPLITT-OUT-R-INt 0 X536-SPLITT-OUT-R-IN 0 z0=5 td=10.0ps
X536 X508-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-IN X536-LSmitll_SPLITT-OUT-X134-LSmitll_DFFT-INt X536-SPLITT-OUT-R-INt LSmitll_SPLITT

t1730 X537-LSmitll_SPLITT-OUT-X135-LSmitll_DFFT-INt 0 X537-LSmitll_SPLITT-OUT-X135-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1731 X537-SPLITT-OUT-R-INt 0 X537-SPLITT-OUT-R-IN 0 z0=5 td=9.8ps
X537 X501-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-IN X537-LSmitll_SPLITT-OUT-X135-LSmitll_DFFT-INt X537-SPLITT-OUT-R-INt LSmitll_SPLITT

t1732 X538-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-INt 0 X538-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1733 X538-SPLITT-OUT-R-INt 0 X538-SPLITT-OUT-R-IN 0 z0=5 td=9.8ps
X538 X462-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-IN X538-LSmitll_SPLITT-OUT-X136-LSmitll_DFFT-INt X538-SPLITT-OUT-R-INt LSmitll_SPLITT

t1734 X539-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-INt 0 X539-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1735 X539-SPLITT-OUT-R-INt 0 X539-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X539 X435-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-IN X539-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-INt X539-SPLITT-OUT-R-INt LSmitll_SPLITT

t1736 X540-LSmitll_SPLITT-OUT-X143-LSmitll_XORT-INt 0 X540-LSmitll_SPLITT-OUT-X143-LSmitll_XORT-IN 0 z0=5 td=0.8ps
t1737 X540-SPLITT-OUT-R-INt 0 X540-SPLITT-OUT-R-IN 0 z0=5 td=9.7ps
X540 X379-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-IN X540-LSmitll_SPLITT-OUT-X143-LSmitll_XORT-INt X540-SPLITT-OUT-R-INt LSmitll_SPLITT

t1738 X541-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-INt 0 X541-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-IN 0 z0=5 td=0.9ps
t1739 X541-SPLITT-OUT-R-INt 0 X541-SPLITT-OUT-R-IN 0 z0=5 td=10.5ps
X541 X382-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-IN X541-LSmitll_SPLITT-OUT-X159-LSmitll_XORT-INt X541-SPLITT-OUT-R-INt LSmitll_SPLITT

t1740 X542-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-INt 0 X542-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-IN 0 z0=5 td=0.4ps
t1741 X542-SPLITT-OUT-R-INt 0 X542-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X542 X366-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-IN X542-LSmitll_SPLITT-OUT-X185-LSmitll_AND2T-INt X542-SPLITT-OUT-R-INt LSmitll_SPLITT

t1742 X543-LSmitll_SPLITT-OUT-X190-LSmitll_AND2T-INt 0 X543-LSmitll_SPLITT-OUT-X190-LSmitll_AND2T-IN 0 z0=5 td=0.7ps
t1743 X543-SPLITT-OUT-R-INt 0 X543-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X543 X486-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-IN X543-LSmitll_SPLITT-OUT-X190-LSmitll_AND2T-INt X543-SPLITT-OUT-R-INt LSmitll_SPLITT

t1744 X544-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-INt 0 X544-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-IN 0 z0=5 td=0.7ps
t1745 X544-SPLITT-OUT-R-INt 0 X544-SPLITT-OUT-R-IN 0 z0=5 td=9.8ps
X544 X372-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-IN X544-LSmitll_SPLITT-OUT-X202-LSmitll_OR2T-INt X544-SPLITT-OUT-R-INt LSmitll_SPLITT

t1746 X545-LSmitll_SPLITT-OUT-X206-LSmitll_OR2T-INt 0 X545-LSmitll_SPLITT-OUT-X206-LSmitll_OR2T-IN 0 z0=5 td=1.0ps
t1747 X545-SPLITT-OUT-R-INt 0 X545-SPLITT-OUT-R-IN 0 z0=5 td=9.9ps
X545 X397-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-IN X545-LSmitll_SPLITT-OUT-X206-LSmitll_OR2T-INt X545-SPLITT-OUT-R-INt LSmitll_SPLITT

t1748 X546-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-INt 0 X546-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1749 X546-SPLITT-OUT-R-INt 0 X546-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X546 X327-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-IN X546-LSmitll_SPLITT-OUT-X225-LSmitll_DFFT-INt X546-SPLITT-OUT-R-INt LSmitll_SPLITT

t1750 X547-LSmitll_SPLITT-OUT-X236-LSmitll_DFFT-INt 0 X547-LSmitll_SPLITT-OUT-X236-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1751 X547-SPLITT-OUT-R-INt 0 X547-SPLITT-OUT-R-IN 0 z0=5 td=10.0ps
X547 X392-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-IN X547-LSmitll_SPLITT-OUT-X236-LSmitll_DFFT-INt X547-SPLITT-OUT-R-INt LSmitll_SPLITT

t1752 X548-LSmitll_SPLITT-OUT-X243-LSmitll_DFFT-INt 0 X548-LSmitll_SPLITT-OUT-X243-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1753 X548-SPLITT-OUT-R-INt 0 X548-SPLITT-OUT-R-IN 0 z0=5 td=9.7ps
X548 X460-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-IN X548-LSmitll_SPLITT-OUT-X243-LSmitll_DFFT-INt X548-SPLITT-OUT-R-INt LSmitll_SPLITT

t1754 X549-LSmitll_SPLITT-OUT-X244-LSmitll_OR2T-INt 0 X549-LSmitll_SPLITT-OUT-X244-LSmitll_OR2T-IN 0 z0=5 td=0.7ps
t1755 X549-SPLITT-OUT-R-INt 0 X549-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X549 X332-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-IN X549-LSmitll_SPLITT-OUT-X244-LSmitll_OR2T-INt X549-SPLITT-OUT-R-INt LSmitll_SPLITT

t1756 X550-LSmitll_SPLITT-OUT-X251-LSmitll_DFFT-INt 0 X550-LSmitll_SPLITT-OUT-X251-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1757 X550-SPLITT-OUT-R-INt 0 X550-SPLITT-OUT-R-IN 0 z0=5 td=10.0ps
X550 X474-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-IN X550-LSmitll_SPLITT-OUT-X251-LSmitll_DFFT-INt X550-SPLITT-OUT-R-INt LSmitll_SPLITT

t1758 X551-LSmitll_SPLITT-OUT-X263-LSmitll_DFFT-INt 0 X551-LSmitll_SPLITT-OUT-X263-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1759 X551-SPLITT-OUT-R-INt 0 X551-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X551 X355-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-IN X551-LSmitll_SPLITT-OUT-X263-LSmitll_DFFT-INt X551-SPLITT-OUT-R-INt LSmitll_SPLITT

t1760 X552-LSmitll_SPLITT-OUT-X265-LSmitll_DFFT-INt 0 X552-LSmitll_SPLITT-OUT-X265-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1761 X552-SPLITT-OUT-R-INt 0 X552-SPLITT-OUT-R-IN 0 z0=5 td=10.1ps
X552 X357-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-IN X552-LSmitll_SPLITT-OUT-X265-LSmitll_DFFT-INt X552-SPLITT-OUT-R-INt LSmitll_SPLITT

t1762 X553-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-INt 0 X553-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
t1763 X553-SPLITT-OUT-R-INt 0 X553-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X553 X352-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-IN X553-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-INt X553-SPLITT-OUT-R-INt LSmitll_SPLITT

t1764 X554-LSmitll_SPLITT-OUT-X281-LSmitll_DFFT-INt 0 X554-LSmitll_SPLITT-OUT-X281-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1765 X554-SPLITT-OUT-R-INt 0 X554-SPLITT-OUT-R-IN 0 z0=5 td=10.1ps
X554 X437-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-IN X554-LSmitll_SPLITT-OUT-X281-LSmitll_DFFT-INt X554-SPLITT-OUT-R-INt LSmitll_SPLITT

t1766 X555-LSmitll_SPLITT-OUT-X286-LSmitll_DFFT-INt 0 X555-LSmitll_SPLITT-OUT-X286-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
t1767 X555-SPLITT-OUT-R-INt 0 X555-SPLITT-OUT-R-IN 0 z0=5 td=9.9ps
X555 X471-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-IN X555-LSmitll_SPLITT-OUT-X286-LSmitll_DFFT-INt X555-SPLITT-OUT-R-INt LSmitll_SPLITT

t1768 X556-LSmitll_SPLITT-OUT-X290-LSmitll_XORT-INt 0 X556-LSmitll_SPLITT-OUT-X290-LSmitll_XORT-IN 0 z0=5 td=0.6ps
t1769 X556-SPLITT-OUT-R-INt 0 X556-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X556 X432-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-IN X556-LSmitll_SPLITT-OUT-X290-LSmitll_XORT-INt X556-SPLITT-OUT-R-INt LSmitll_SPLITT

t1770 X557-LSmitll_SPLITT-OUT-X292-LSmitll_OR2T-INt 0 X557-LSmitll_SPLITT-OUT-X292-LSmitll_OR2T-IN 0 z0=5 td=0.9ps
t1771 X557-SPLITT-OUT-R-INt 0 X557-SPLITT-OUT-R-IN 0 z0=5 td=10.5ps
X557 X395-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-IN X557-LSmitll_SPLITT-OUT-X292-LSmitll_OR2T-INt X557-SPLITT-OUT-R-INt LSmitll_SPLITT

t1772 X558-LSmitll_SPLITT-OUT-X293-LSmitll_DFFT-INt 0 X558-LSmitll_SPLITT-OUT-X293-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1773 X558-SPLITT-OUT-R-INt 0 X558-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X558 X457-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-IN X558-LSmitll_SPLITT-OUT-X293-LSmitll_DFFT-INt X558-SPLITT-OUT-R-INt LSmitll_SPLITT

t1774 X559-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-INt 0 X559-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1775 X559-SPLITT-OUT-R-INt 0 X559-SPLITT-OUT-R-IN 0 z0=5 td=10.2ps
X559 X445-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-IN X559-LSmitll_SPLITT-OUT-X297-LSmitll_DFFT-INt X559-SPLITT-OUT-R-INt LSmitll_SPLITT

t1776 X560-LSmitll_SPLITT-OUT-X299-LSmitll_DFFT-INt 0 X560-LSmitll_SPLITT-OUT-X299-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
t1777 X560-SPLITT-OUT-R-INt 0 X560-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X560 X419-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-IN X560-LSmitll_SPLITT-OUT-X299-LSmitll_DFFT-INt X560-SPLITT-OUT-R-INt LSmitll_SPLITT

t1778 X561-LSmitll_SPLITT-OUT-X302-LSmitll_DFFT-INt 0 X561-LSmitll_SPLITT-OUT-X302-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1779 X561-SPLITT-OUT-R-INt 0 X561-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X561 X496-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-IN X561-LSmitll_SPLITT-OUT-X302-LSmitll_DFFT-INt X561-SPLITT-OUT-R-INt LSmitll_SPLITT

t1780 X562-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-INt 0 X562-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1781 X562-SPLITT-OUT-R-INt 0 X562-SPLITT-OUT-R-IN 0 z0=5 td=9.8ps
X562 X425-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-IN X562-LSmitll_SPLITT-OUT-X304-LSmitll_DFFT-INt X562-SPLITT-OUT-R-INt LSmitll_SPLITT

t1782 X563-LSmitll_SPLITT-OUT-X307-LSmitll_DFFT-INt 0 X563-LSmitll_SPLITT-OUT-X307-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1783 X563-SPLITT-OUT-R-INt 0 X563-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X563 X499-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-IN X563-LSmitll_SPLITT-OUT-X307-LSmitll_DFFT-INt X563-SPLITT-OUT-R-INt LSmitll_SPLITT

t1784 X564-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-INt 0 X564-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-IN 0 z0=5 td=10.7ps
t1785 X564-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-INt 0 X564-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-IN 0 z0=5 td=11.7ps
X564 GCLK X564-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-INt X564-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-INt LSmitll_SPLITT

* PTLs from input pads
t868 GCLKt 0 GCLK 0 z0=5 td=13.3ps

t568 Imm3t 0 Imm3 0 z0=5 td=5.8ps
t572 Imm2t 0 Imm2 0 z0=5 td=11.6ps
t576 Imm1t 0 Imm1 0 z0=5 td=14.7ps
t580 Imm0t 0 Imm0 0 z0=5 td=8.0ps
t584 select1t 0 select1 0 z0=5 td=5.6ps
t588 select0t 0 select0 0 z0=5 td=6.7ps
t604 addr1t 0 addr1 0 z0=5 td=8.2ps
t592 addr0t 0 addr0 0 z0=5 td=7.4ps
t596 readt 0 read 0 z0=5 td=10.5ps
t600 write_flagst 0 write_flags 0 z0=5 td=10.3ps

t616 Op_Aritht 0 Op_Arith 0 z0=5 td=6.1ps
t628 Op_Andt 0 Op_And 0 z0=5 td=2.6ps
t624 Op_Xort 0 Op_Xor 0 z0=5 td=6.6ps
t612 Cmpl_b1t 0 Cmpl_b1 0 z0=5 td=11.8ps
t608 Cmpl_b0t 0 Cmpl_b0 0 z0=5 td=15.1ps
t620 Cint 0 Cin 0 z0=5 td=9.3ps

* PTLs to output pads
t1042 reg1_out3_padt 0 reg1_out3_pad 0 z0=5 td=4.4ps
t1040 reg1_out2_padt 0 reg1_out2_pad 0 z0=5 td=3.3ps
t1038 reg1_out1_padt 0 reg1_out1_pad 0 z0=5 td=7.7ps
t1036 reg1_out0_padt 0 reg1_out0_pad 0 z0=5 td=8.4ps

t1050 reg2_out3_padt 0 reg2_out3_pad 0 z0=5 td=3.2ps
t1048 reg2_out2_padt 0 reg2_out2_pad 0 z0=5 td=3.9ps
t1046 reg2_out1_padt 0 reg2_out1_pad 0 z0=5 td=11.1ps
t1044 reg2_out0_padt 0 reg2_out0_pad 0 z0=5 td=3.4ps

t1056 regFlags_out2_padt 0 regFlags_out2_pad 0 z0=5 td=5.3ps
t1053 regFlags_out1_padt 0 regFlags_out1_pad 0 z0=5 td=2.6ps
t1052 regFlags_out0_padt 0 regFlags_out0_pad 0 z0=5 td=3.5ps

t1055 regFlags_out2t 0 regFlags_out2 0 z0=5 td=10.4ps
t1054 regFlags_out1t 0 regFlags_out1 0 z0=5 td=6.8ps
t1051 regFlags_out0t 0 regFlags_out0 0 z0=5 td=2.4ps

.ends ALU_Reg_file_final_route