* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

* The cell is not designed to be connected directly to passive transmission lines

*$Ports  a b clk q
.subckt LSMITLL_AND2 a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=2.01
.param B3=1.91
.param B4=1.26
.param B5=1.57
.param B6=1.19
.param B7=B1
.param B8=B2
.param B9=B3
.param B10=B4
.param B11=B5
.param B12=B6
.param B13=IC
.param B14=2.06
.param B15=IC

.param IB1=BiasCoef*Ic0*B1
.param IB2=123u
.param IB3=IB1
.param IB4=IB2
.param IB5=BiasCoef*Ic0*B13
.param IB6=133u
.param IB7=BiasCoef*Ic0*B15

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB

.param L1=Phi0/(4*IC*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(B3*Ic0)
.param L4=1p
.param L5=Phi0/(2*B5*Ic0)
.param L6=L1
.param L7=L2
.param L8=L3
.param L9=L4
.param L10=L5
.param L11=Phi0/(4*IC*Ic0)
.param L12=Phi0/(2*B13*Ic0)
.param L13=1p
.param L14=1p
.param L15=Phi0/(4*IC*Ic0)

.param LP1=LP
.param LP3=LP
.param LP5=LP
.param LP7=LP
.param LP9=LP
.param LP11=LP
.param LP13=LP
.param LP14=LP
.param LP15=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet
.param LRB13=(RB13/Rsheet)*Lsheet
.param LRB14=(RB14/Rsheet)*Lsheet
.param LRB15=(RB15/Rsheet)*Lsheet

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 5 6 jjmit area=B3
B4 8 9 jjmit area=B4
B5 8 11 jjmit area=B5
B6 12 13 jjmit area=B6
B7 14 15 jjmit area=B7
B8 17 18 jjmit area=B8
B9 18 19 jjmit area=B9
B10 21 22 jjmit area=B10
B11 21 23 jjmit area=B11
B12 24 13 jjmit area=B12
B13 25 26 jjmit area=B13
B14 31 32 jjmit area=B14
B15 28 29 jjmit area=B15

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 16 pwl(0 0 5p IB3)
IB4 0 20 pwl(0 0 5p IB4)
IB5 0 27 pwl(0 0 5p IB5)
IB6 0 33 pwl(0 0 5p IB6)
IB7 0 30 pwl(0 0 5p IB7)

LB1 3 1 LB1
LB2 7 5 LB2
LB3 16 14 LB3
LB4 20 18 LB4
LB5 27 25 LB5
LB6 30 28 LB6
LB7 33 31 LB7

LP1 2 0 4.864E-13
LP3 6 0 5.474E-13
LP5 11 0 5.279E-13
LP7 15 0 4.901E-13
LP9 19 0 5.414E-13
LP11 23 0 5.306E-13
LP13 26 0 5.084E-13
LP14 32 0 5.329E-13
LP15 29 0 4.92E-13

L1 a 1 2.075E-12
L2 1 4 2.812E-12
L3 5 8 9.756E-12
L4 9 10 1.079E-12
L5 8 12 3.105E-12
L6 b 14 2.073E-12
L7 14 17 2.811E-12
L8 18 21 9.768E-12
L9 22 10 1.084E-12
L10 21 24 3.095E-12
L11 clk 25 2.063E-12
L12 25 31 2.96E-12
L13 31 10 1.002E-12
L14 13 28 1.06E-12
L15 28 q 2.069E-12

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 5 LRB2
RB3 5 105 RB3
LRB3 105 0 LRB3
RB4 8 109 RB4
LRB4 109 9 LRB4
RB5 8 108 RB5
LRB5 108 0 LRB5
RB6 12 112 RB6
LRB6 112 13 LRB6
RB7 14 114 RB7
LRB7 114 0 LRB7
RB8 17 117 RB8
LRB8 117 18 LRB8
RB9 18 118 RB9
LRB9 118 0 LRB9
RB10 21 122 RB10
LRB10 122 22 LRB10
RB11 21 121 RB11
LRB11 121 0 LRB11
RB12 24 124 RB12
LRB12 124 13 LRB12
RB13 25 125 RB13
LRB13 125 0 LRB13
RB14 31 131 RB14
LRB14 131 0 LRB14
RB15 28 128 RB15
LRB15 128 0 LRB15
.ends LSMITLL_AND2


*$Ports		a b clk q
.SUBCKT LSMITLL_OR2 a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7

.param B1=2.5
.param B2=2.22
.param B3=1.86
.param B4=B1
.param B5=B2
.param B6=B3
.param B7=2.28
.param B8=2.09
.param B9=2.5
.param B10=1.52
.param B11=1.60
.param B12=2.5

.param IB1=175u
.param IB2=IB1
.param IB3=304u
.param IB4=142u
.param IB5=175u
.param IB6=175u

.param L1=Phi0/(4*IC*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=1p
.param L4=L1
.param L5=L2
.param L6=L3
.param L7=Phi0/(2*B2*Ic0)
.param L8=Phi0/(B8*Ic0)
.param L9=Phi0/(4*IC*Ic0)
.param L10=Phi0/(2*B9*Ic0)
.param L11=Phi0/(2*B11*Ic0)
.param L12=Phi0/(4*IC*Ic0)

.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10 
.param RB11=B0Rs/B11 
.param RB12=B0Rs/B12 
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP 
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP 
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet+LP
.param LRB12=(RB12/Rsheet)*Lsheet+LP

L1 a 1 2.051E-12
L2 1 4 3.232E-12
L3 4 6 1.198E-12
L4 b 8 2.046E-12 
L5 8 11 3.242E-12
L6 11 13 1.191E-12
L7 7 15 3.341E-12
L8 16 19 7.998E-12
L9 clk 20 2.062E-12
L10 20 23 3.408E-12
L11 19 25 3.54E-12
L12 25 q 2.05E-12

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 6 7 jjmit area=B3
B4 8 9 jjmit area=B4
B5 11 12 jjmit area=B5
B6 13 7 jjmit area=B6
B7 15 16 jjmit area=B7
B8 16 17 jjmit area=B8
B9 20 21 jjmit area=B9
B10 23 19 jjmit area=B10
B11 19 24 jjmit area=B11
B12 25 26 jjmit area=B12

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)
IB3 0 14 pwl(0 0 5p IB3)
IB4 0 18 pwl(0 0 5p IB4)
IB5 0 22 pwl(0 0 5p IB5)
IB6 0 27 pwl(0 0 5p IB6)

LB1 1 3 LB
LB2 8 10 LB
LB3 7 14 LB
LB4 16 18 LB
LB5 20 22 LB
LB6 25 27 LB

LP1 2 0 5.253E-13
LP2 5 0 5.141E-13
LP4 9 0 5.352E-13
LP5 12 0 5.154E-13
LP8 17 0 4.905E-13
LP9 21 0 5.216E-13
LP11 24 0 5.649E-13
LP12 26 0 5.28E-13

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 0 LRB2
RB3 6 105 RB3
LRB3 105 7 LRB3
RB4 8 108 RB4
LRB4 108 0 LRB4
RB5 11 111 RB5
LRB5 111 0 LRB5
RB6 13 113 RB6
LRB6 113 7 LRB6
RB7 15 115 RB7
LRB7 115 16 LRB7
RB8 16 116 RB8
LRB8 116 0 LRB8
RB9 20 120 RB9
LRB9 120 0 LRB9
RB10 23 123 RB10
LRB10 123 19 LRB10
RB11 19 119 RB11
LRB11 119 0 LRB11
RB12 25 125 RB12
LRB12 125 0 LRB12
.ends LSMITLL_OR2


*$Ports a b clk q
.subckt LSmitll_XOR	a	b	clk 	q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.70
.param B1=2.5
.param B2=2.09
.param B3=1.71
.param B4=B1
.param B5=B2
.param B6=B3
.param B7=1.62
.param B8=2.5
.param B9=1.45
.param B10=0.89
.param B11=2.5
.param IB1=175u
.param IB2=112u
.param IB3=IB1
.param IB4=IB2
.param IB5=175u
.param IB6=175u
.param L1=Phi0/(4*IC*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=1.2p
.param L4=Phi0/(B2*Ic0)
.param L5=L1
.param L6=L2
.param L7=L3
.param L8=L4
.param L9=1.2p
.param L10=Phi0/(4*IC*Ic0)
.param L11=Phi0/(2*B8*Ic0)
.param L12=Phi0/(2*B10*Ic0)
.param L13=Phi0/(4*IC*Ic0)
.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3          
.param RB4=B0Rs/B4         
.param RB5=B0Rs/B5         
.param RB6=B0Rs/B6          
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8         
.param RB9=B0Rs/B9         
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet+LP
B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 25 6 jjmit area=B3
B4 9 10 jjmit area=B4
B5 12 13 jjmit area=B5
B6 26 14 jjmit area=B6
B7 27 16 jjmit area=B7
B8 17 18 jjmit area=B8
B9 20 16 jjmit area=B9
B10 16 21 jjmit area=B10
B11 22 23 jjmit area=B11
IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 11 pwl(0 0 5p IB3)
IB4 0 15 pwl(0 0 5p IB4)
IB5 0 19 pwl(0 0 5p IB5)
IB6 0 24 pwl(0 0 5p IB6)
LB1 3 1 LB
LB2 7 6 LB
LB3 11 9 LB
LB4 15 14 LB
LB5 19 17 LB
LB6 24 22 LB
L1 a 1 2.06E-12
L2 1 4 3.233E-12
L3 4 25 1.419E-12
L4 6 8 6.051E-12
L5 b 9 2.092E-12
L6 9 12 3.221E-12
L7 12 26 1.384E-12
L8 14 8 6.059E-12
L9 8 27 1.301E-12
L10 clk 17 2.082E-12
L11 17 20 1.43E-12
L12 16 22 3.892E-12
L13 22 q 2.077E-12
LP1 2 0 5.508E-13
LP2 5 0 4.769E-13
LP4 10 0 4.767E-13
LP5 13 0 4.812E-13
LP8 18 0 4.526E-13
LP10 21 0 5.69E-13
LP11 23 0 4.746E-13
RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 0 LRB2
RB3 4 106 RB3
LRB3 106 6 LRB3
RB4 9 109 RB4
LRB4 109 0 LRB4
RB5 12 112 RB5
LRB5 112 0 LRB5
RB6 12 114 RB6
LRB6 114 14 LRB6
RB7 8 108 RB7
LRB7 108 16 LRB7
RB8 17 117 RB8
LRB8 117 0 LRB8
RB9 20 120 RB9
LRB9 120 16 LRB9
RB10 16 116 RB10
LRB10 116 0 LRB10
RB11 22 122 RB11
LRB11 122 0 LRB11
.ends LSmitll_XOR


*$Ports  a clk q
.subckt LSMITLL_NOT a clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=2.57
.param B3=1.07
.param B4=IC
.param B5=1.34
.param B6=3.03
.param B7=1.38
.param B8=0.8
.param B9=IC

.param IB1=BiasCoef*Ic0*B1
.param IB2=87u
.param IB3=257u
.param IB4=BiasCoef*Ic0*B4
.param IB5=BiasCoef*Ic0*B9

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9

.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet

.param RD=4
.param LRD=2p

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 7 8 jjmit area=B3
B4 13 14 jjmit area=B4
B5 17 18 jjmit area=B5
B6 10 11 jjmit area=B6
B7 20 18 jjmit area=B7
B8 18 19 jjmit area=B8
B9 21 22 jjmit area=B9

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 9 pwl(0 0 5p IB3)
IB4 0 15 pwl(0 0 5p IB4)
IB5 0 23 pwl(0 0 5p IB5)

LB1 3 1 LB1
LB2 6 4 LB2
LB3 8 9 LB3
LB4 13 15 LB4
LB5 21 23 LB5

L1 a 1 2.062E-12
L2 1 4 1.889E-12
L3 4 7 2.72E-12
L4 clk 13 2.057E-12
L5 13 16 1.029E-12
L6 16 17 1.241E-12
L7 16 12 1.973E-12
L8 10 12 1.003E-12
L9 10 8 7.524E-12
L10 8 20 1.234E-12
L11 18 21 2.607E-12
L12 21 q 2.062E-12

LP1 2 0 5.271E-13
LP2 5 0 5.237E-13
LP4 14 0 4.759E-13
LP6 11 0 5.021E-13
LP8 19 0 6.33E-13
LP9 22 0 4.749E-13

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 5 LRB2
RB3 7 107 RB3
LRB3 107 8 LRB3
RB4 13 113 RB4
LRB4 113 0 LRB4
RB5 17 117 RB5
LRB5 117 18 LRB5
RB6 10 110 RB6
LRB6 110 0 LRB6
RB7 20 120 RB7
LRB7 120 18 LRB7
RB8 18 118 RB8
LRB8 118 0 LRB8
RB9 21 121 RB9
LRB9 121 0 LRB9
LRD 12 112 LRD
RD 112 0 RD
.ends LSMITLL_NOT


*$Ports a q0 q1
.subckt LSmitll_SPLIT a q0 q1
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7
.param RD=1.36

.param B1=2.5
.param B2=3.0
.param B3=2.5
.param B4=2.5

.param IB1=175u
.param IB2=280u
.param IB3=175u
.param IB4=175u

.param L1=Lptl
.param L2=Phi0/(2*B1*Ic0)
.param L3=(Phi0/(2*B2*Ic0))/2
.param L4=L3
.param L5=Lptl
.param L6=L3
.param L7=Lptl

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 10 pwl(0 0 5p IB3)
IB4 0 13 pwl(0 0 5p IB4)
LB1 3 1 9.175E-13
LB2 6 4 7.666E-13
LB3 10 8 1.928E-12
LB4 13 11 8.786E-13

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 8 9 jjmit area=B3
B4 11 12 jjmit area=B4
L1 a 1 2.063E-12
L2 1 4 3.637E-12
L3 4 7 1.278E-12
L4 7 8 1.305E-12
L5 8 q0 2.05E-12
L6 7 11 1.315E-12
L7 11 q1 2.06E-12

LP1 2 0 4.676E-13
LP2 5 0 4.498E-13
LP3 9 0 5.183E-13
LP4 12 0 4.639E-13
RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 0 LRB2
RB3 8 108 RB3
LRB3 108 0 LRB3
RB4 11 111 RB4
LRB4 111 0 LRB4
.ends LSmitll_SPLIT


*$Ports a q
.subckt LSMITLL_BUFF a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC
.param B3=IC
.param B4=IC
.param IB1=B1*Ic0*BiasCoef
.param IB2=B2*Ic0*0.95
.param IB3=B3*Ic0*0.95
.param IB4=B4*Ic0*BiasCoef
.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param L1=Phi0/(4*IC*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(2*B2*Ic0)
.param L4=Phi0/(2*B3*Ic0)
.param L5=Phi0/(4*IC*Ic0)
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP
.param LP3=LP
.param LP4=LP

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 7 8 jjmit area=B3
B4 10 11 jjmit area=B4

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 9 pwl(0 0 5p IB3)
IB4 0 12 pwl(0 0 5p IB4)

L1 a 1 2.057E-12
L2 1 4 4.026E-12
L3 4 7 4.155E-12
L4 7 10 4.057E-12
L5 10 q 2.057E-12

LP1 2 0 5.283E-13
LP2 5 0 5.327E-13
LP3 8 0 5.084E-13
LP4 11 0 5.269E-13

LB1 1 3 LB1
LB2 4 6 LB2
LB3 7 9 LB3
LB4 10 12 LB4

RB1 1 101 RB1
RB2 4 104 RB2
RB3 7 107 RB3
RB4 10 110 RB4

LRB1 101 0 LRB1
LRB2 104 0 LRB2
LRB3 107 0 LRB3
LRB4 110 0 LRB4
.ends LSMITLL_BUFF


*$Ports		a		clk		q
.subckt LSmitll_DFF	  a	clk q	
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.70

.param B1=2.5
.param B2=1.61
.param B3=1.54
.param B4=1.69
.param B5=1.38
.param B6=2.5
.param B7=2.5

.param IB1=175u     
.param IB2=173u      
.param IB3=175u            
.param IB4=175u        

.param L1=Phi0/(4*IC*Ic0)               
.param L2=Phi0/(2*B1*Ic0)         
.param L3=Phi0/(B3*Ic0)       
.param L4=Phi0/(2*B6*Ic0)      
.param L5=Phi0/(4*IC*Ic0)     
.param L6=Phi0/(2*B4*Ic0)       
.param L7=Phi0/(4*B7*Ic0)         
.param LB1=LB            
.param LB2=LB           
.param LB3=LB           
.param LB4=LB        
.param LP1=LP         
.param LP3=LP          
.param LP4=LP         
.param LP6=LP          
.param LP7=LP          
.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3          
.param RB4=B0Rs/B4         
.param RB5=B0Rs/B5         
.param RB6=B0Rs/B6          
.param RB7=B0Rs/B7
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 5 6 jjmit area=B3
B4 8 9 jjmit area=B4
B5 10 8 jjmit area=B5
B6 11 12 jjmit area=B6
B7 14 15 jjmit area=B7

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 13 pwl(0 0 5p IB3)
IB4 0 16 pwl(0 0 5p IB4)

LB1 3 1 LB1
LB2 7 5 LB2
LB3 11 13 LB3
LB4 16 14 LB4

L1 a 1 2.059E-12
L2 1 4 4.123E-12
L3 5 8 6.873E-12
L4 10 11 5.195E-12
L5 clk 11 2.071E-12
L6 8 14 3.287E-12
L7 14 q 2.066E-12

LP1 2 0 5.042E-13    
LP3 6 0 5.799E-13    
LP4 9 0 5.733E-13    
LP6 12 0 4.605E-13    
LP7 15 0 4.961E-13    

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 5 LRB2
RB3 5 105 RB3
LRB3 105 0 LRB3
RB4 8 108 RB4
LRB4 108 0 LRB4
RB5 10 110 RB5
LRB5 110 8 LRB5
RB6 11 111 RB6
LRB6 111 0 LRB6
RB7 14 114 RB7
LRB7 114 0 LRB7
.ends LSmitll_DFF

*$Ports 		 q
.subckt LSMITLL_Always0_async_noA  q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7
.param B1=IC
.param IB1=B1*Ic0*BiasCoef
.param L1=Phi0/(2*B1*Ic0)
.param L2=Phi0/(4*B1*Ic0)
.param LB1=LB
.param RB1=B0Rs/B1   
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LP1=LP
.param R1=2

B1 2 3 jjmit area=B1
IB1 0 5 pwl(0 0 5p IB1)
L1 1 2 1.397E-12
L2 2 q 2.465E-12
R1 1 0 R1
LB1 2 4 3.177E-12
LP1 3 0 5.306E-13
RB1 2 102 RB1
LRB1 102 0 LRB1
.ends LSMITLL_Always0_async_noA

*$Ports 			a q
.subckt LSMITLL_Always0_async a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7
.param B1=IC
.param B2=IC
.param IB1=B1*Ic0*BiasCoef
.param IB2=B2*Ic0*BiasCoef
.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(2*B2*Ic0)
.param L4=Phi0/(4*B2*Ic0)
.param LB1=LB
.param LB2=LB
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP
.param R1=2
.param R2=2

B1 1 2 jjmit area=B1
B2 6 7 jjmit area=B2
IB1 0 3 pwl(0 0 5p IB1)
IB2 0 8 pwl(0 0 5p IB2)
L1 a 1 2.47E-12
L2 1 4 1.4E-12
L3 5 6 2.948E-12
L4 6 q 3.768E-12
R1 4 0 R1
R2 5 0 R2
LB1 1 3 2.199E-12
LB2 6 8 1.087E-12
LP1 2 0 5.282E-13
LP2 7 0 4.908E-13
RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 6 106 RB2
LRB2 106 0 LRB2
.ends LSMITLL_Always0_async


*$Ports 			clk q
.subckt LSMITLL_Always0_sync_noA clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7
.param B1=IC
.param B2=IC
.param IB1=B1*Ic0*BiasCoef
.param IB2=B2*Ic0*BiasCoef
.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(2*B2*Ic0)
.param L4=Phi0/(4*B2*Ic0)
.param LB1=LB
.param LB2=LB
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP
.param R1=2
.param R2=2

B1 1 2 jjmit area=B1
B2 6 7 jjmit area=B2
IB1 0 3 pwl(0 0 5p IB1)
IB2 0 8 pwl(0 0 5p IB2)
L1 clk 1 2.507E-12
L2 1 4 1.057E-12
L3 5 6 1.062E-12
L4 6 q 3.747E-12
R1 4 0 R1
R2 5 0 R2
LB1 1 3 2.133E-12
LB2 6 8 2.17E-12
LP1 2 0 4.927E-13
LP2 7 0 4.925E-13
RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 6 106 RB2
LRB2 106 0 LRB2
.ends LSMITLL_Always0_sync_noA

*$Ports 			a clk q
.subckt LSMITLL_Always0_sync a clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7
.param B1=IC
.param B2=IC
.param B3=IC
.param IB1=B1*Ic0*BiasCoef
.param IB2=B2*Ic0*BiasCoef
.param IB3=B3*Ic0*BiasCoef
.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(4*B2*Ic0)
.param L4=Phi0/(2*B2*Ic0)
.param L5=Phi0/(2*B3*Ic0)
.param L6=Phi0/(4*B3*Ic0)
.param LB1=LB
.param LB2=LB
.param LB3=LB
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP
.param LP3=LP
.param R1=2
.param R2=2
.param R3=2

B1 1 2 jjmit area=B1
B2 5 6 jjmit area=B2
B3 10 11 jjmit area=B3
IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 12 pwl(0 0 5p IB3)
L1 a 1 3.78E-12
L2 1 4 1.016E-12
L3 clk 5 2.5E-12
L4 5 8 1.048E-12
L5 9 10 1.005E-12
L6 10 q 2.488E-12
R1 4 0 R1
R2 8 0 R2
R3 9 0 R3
LB1 1 3 1.243E-12
LB2 5 7 2.181E-12
LB3 10 12 5.092E-12
LP1 2 0 4.931E-13
LP2 6 0 4.919E-13
LP3 11 0 5.015E-13
RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 5 105 RB2
LRB2 105 0 LRB2
RB3 10 110 RB3
LRB3 110 0 LRB3
.ends LSMITLL_Always0_sync


*$Ports a b clk q
.subckt LSmitll_NDRO a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=2.5
.param B2=1.99
.param B3=2.2
.param B4=2.5
.param B5=2.35
.param B6=3.24
.param B7=0.74
.param B8=2.5
.param B9=1.17
.param B10=1.09
.param B11=2.5

.param IB1=175u
.param IB2=271u
.param IB3=175u
.param IB4=175u
.param IB5=136u
.param IB6=175u

.param L1=Phi0/(4*IC*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(2*B3*Ic0)
.param L4=Phi0/(4*IC*Ic0)
.param L5=Phi0/(2*B4*Ic0)
.param L6=Phi0/(2*B6*Ic0)
.param L7=1p
.param L8=1p
.param L9=Phi0/(4*IC*Ic0)
.param L10=Phi0/(2*B8*Ic0)
.param L11=Phi0/(2*B10*Ic0)
.param L12=Phi0/(4*IC*Ic0)

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet+LP

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB

B1 1 2 jjmit area=B1
B2 3 4 jjmit area=B2
B3 4 5 jjmit area=B3
B4 7 8 jjmit area=B4
B5 9 10 jjmit area=B5
B6 10 11 jjmit area=B6
B7 6 12 jjmit area=B7
B8 14 15 jjmit area=B8
B9 14 16 jjmit area=B9
B10 17 18 jjmit area=B10
B11 19 20 jjmit area=B11

IB1 0 21 pwl(0 0 5p IB1)
IB2 0 22 pwl(0 0 5p IB2)
IB3 0 23 pwl(0 0 5p IB3)
IB4 0 24 pwl(0 0 5p IB4)
IB5 0 25 pwl(0 0 5p IB5)
IB6 0 26 pwl(0 0 5p IB6)

LB1 1 21 LB1
LB2 4 22 LB2
LB3 7 23 LB3
LB4 14 24 LB4
LB5 13 25 LB5
LB6 19 26 LB6

L1 a 1 2.067E-12
L2 1 3 9.786E-13
L3 4 6 2.693E-12
L4 b 7 2.068E-12
L5 7 9 2.319E-12
L6 10 6 3.438E-12
L7 12 13 1.12E-12
L8 13 17 1.028E-12
L9 clk 14 2.106E-12
L10 16 17 3.135E-12
L11 17 19 3.223E-12
L12 19 q 2.071E-12

LP1 2 0 5.174E-13
LP3 5 0 5.135E-13
LP4 8 0 4.756E-13
LP6 11 0 4.841E-13
LP8 15 0 4.705E-13
LP10 18 0 5.961E-13
LP11 20 0 4.832E-13

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 3 103 RB2
LRB2 103 4 LRB2
RB3 4 104 RB3
LRB3 104 0 LRB3
RB4 7 107 RB4
LRB4 107 0 LRB4
RB5 9 109 RB5
LRB5 109 10 LRB5
RB6 10 110 RB6
LRB6 110 0 LRB6
RB7 6 106 RB7
LRB7 106 12 LRB7
RB8 14 114 RB8
LRB8 114 0 LRB8
RB9 14 116 RB9
LRB9 116 16 LRB9
RB10 17 117 RB10
LRB10 117 0 LRB10
RB11 19 119 RB11
LRB11 119 0 LRB11
.ends LSmitll_NDRO


*$Ports				   a b q
.subckt LSmitll_MERGE a b q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.70
.param RD=1.36

.param B1=IC
.param B2=2.5
.param B3=1.92
.param B4=B1
.param B5=B2
.param B6=B3
.param B7=2.53
.param B8=IC

.param IB1=BiasCoef*Ic0*B1
.param IB2=IB1
.param IB3=254E-6
.param IB4=192E-6
.param IB5=BiasCoef*Ic0*B8

.param L1=Phi0/(4*IC*Ic0)
.param L2=3.173E-12
.param L3=1.2E-12
.param L4=L1
.param L5=L2
.param L6=L3
.param L7=5.354E-12
.param L8=4.456E-12
.param L9=Phi0/(4*B8*Ic0)

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB

.param LP1=LP
.param LP2=LP
.param LP4=LP
.param LP5=LP
.param LP7=LP
.param LP8=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 4 6 jjmit area=B3
B4 8 9 jjmit area=B4
B5 11 12 jjmit area=B5
B6 11 13 jjmit area=B6
B7 15 16 jjmit area=B7
B8 18 19 jjmit area=B8

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)
IB3 0 14 pwl(0 0 5p IB3)
IB4 0 17 pwl(0 0 5p IB4)
IB5 0 20 pwl(0 0 5p IB5)

L1 a 1 2.117E-12
L2 1 4 3.17E-12
L3 6 7 1.234E-12
L4 b 8 2.082E-12
L5 8 11 3.165E-12
L6 13 7 1.224E-12
L7 7 15 5.299E-12
L8 15 18 4.489E-12
L9 18 q 2.077E-12

LP1 2 0 4.652E-13
LP2 5 0 4.457E-13
LP4 9 0 5.293E-13
LP5 12 0 4.452E-13
LP7 16 0 5.039E-13
LP8 19 0 4.984E-13

LB1 1 3 LB1
LB2 8 10 LB2
LB3 7 14 LB3
LB4 15 17 LB4
LB5 18 20 LB5

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 0 LRB2
RB3 4 106 RB3
LRB3 106 6 LRB3
RB4 8 108 RB4
LRB4 108 0 LRB4
RB5 11 111 RB5
LRB5 111 0 LRB5
RB6 11 113 RB6
LRB6 113 13 LRB6
RB7 15 115 RB7
LRB7 115 0 LRB7
RB8 18 118 RB8
LRB8 118 0 LRB8
.ends LSmitll_MERGE

*$Ports  a b clk q
.subckt LSMITLL_XNOR a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7

.param B1=2.5
.param B2=2.66
.param B3=2.34
.param B4=B1
.param B5=B2
.param B6=B3
.param B7=2.31
.param B8=3.15
.param B9=2.5
.param B10=2.58
.param B11=1.44
.param B12=2.60
.param B13=2.71
.param B14=1.63
.param B15=0.95
.param B16=1.44
.param B17=1.40
.param B18=2.5

.param IB1=175E-6
.param IB2=153E-6
.param IB3=IB1
.param IB4=IB2
.param IB5=175E-6
.param IB6=260E-6
.param IB7=56E-6
.param IB8=248E-6
.param IB9=51E-6
.param IB10=175E-6

.param L1=Lptl
.param L2=Phi0/(2*B1*Ic0)
.param L3=1p
.param L4=Phi0/(B2*Ic0)
.param L5=L1
.param L6=L2
.param L7=L3
.param L8=L4
.param L9=1p
.param L10=Lptl
.param L11=Phi0/(2*B9*Ic0)
.param L12=1p
.param L13=1p
.param L14=Phi0/(2*B10*Ic0)
.param L15=Phi0/(4*B12*Ic0)
.param L16=Phi0/(4*B12*Ic0)
.param L17=Phi0/(B13*Ic0)
.param L18=1p
.param L20=1p
.param L21=0.5p
.param L22=Phi0/(B16*Ic0)
.param L23=Phi0/(4*B16*Ic0)
.param L24=Phi0/(2*B17*Ic0)
.param L25=Lptl

.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3          
.param RB4=B0Rs/B4         
.param RB5=B0Rs/B5         
.param RB6=B0Rs/B6          
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8         
.param RB9=B0Rs/B9         
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15
.param RB16=B0Rs/B16
.param RB17=B0Rs/B17
.param RB18=B0Rs/B18
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet
.param LRB13=(RB13/Rsheet)*Lsheet
.param LRB14=(RB14/Rsheet)*Lsheet
.param LRB15=(RB15/Rsheet)*Lsheet
.param LRB16=(RB16/Rsheet)*Lsheet
.param LRB17=(RB17/Rsheet)*Lsheet
.param LRB18=(RB18/Rsheet)*Lsheet

B1 1 2 jjmit area=B1
B2 3 4 jjmit area=B2
B3 5 6 jjmit area=B3
B4 8 9 jjmit area=B4
B5 10 11 jjmit area=B5
B6 12 13 jjmit area=B6
B7 14 15 jjmit area=B7
B8 15 16 jjmit area=B8
B9 17 18 jjmit area=B9
B10 19 20 jjmit area=B10
B11 22 15 jjmit area=B11
B12 23 24 jjmit area=B12
B13 26 27 jjmit area=B13
B14 29 34 jjmit area=B14
B15 34 31 jjmit area=B15
B16 28 33 jjmit area=B16
B17 35 36 jjmit area=B17
B18 37 38 jjmit area=B18

LP1 2 0 5.29E-13
LP2 4 0 4.956E-13
LP4 9 0 4.424E-13
LP5 11 0 5.101E-13
LP8 16 0 5.051E-13
LP9 18 0 5.321E-13
LP10 20 0 5.07E-13
LP12 24 0 5.287E-13
LP13 27 0 5.393E-13
LP17 36 0 5.753E-13
LP18 38 0 5.361E-13

IB1 0 1 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 8 pwl(0 0 5p IB3)
IB4 0 13 pwl(0 0 5p IB4)
IB5 0 17 pwl(0 0 5p IB5)
IB6 0 19 pwl(0 0 5p IB6)
IB7 0 25 pwl(0 0 5p IB7)
IB8 0 34 pwl(0 0 5p IB8)
IB9 0 35 pwl(0 0 5p IB9)
IB10 0 37 pwl(0 0 5p IB10)

L1 a 1 2.058E-12
L2 1 3 2.395E-12
L3 3 5 1.108E-12
L4 6 7 4.1E-12
L5 b 8 2.104E-12
L6 8 10 2.374E-12
L7 10 12 9.887E-13
L8 13 7 4.048E-12
L9 7 14 1.15E-12
L10 clk 17 2.041E-12
L11 17 19 3.442E-12
L12 19 21 8.703E-13
L13 21 22 1.117E-12
L14 21 23 2.107E-12
L15 23 25 1.641E-12
L16 25 26 1.335E-12
L17 26 28 5.203E-12
L18 15 29 1.494E-12
L20 31 32 2.081E-12
L21 33 32 9.13E-13
L22 34 28 6.448E-12
L23 32 35 1.012E-12
L24 35 37 3.546E-12
L25 37 q 2.034E-12

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 3 103 RB2
LRB2 103 0 LRB2
RB3 5 105 RB3
LRB3 105 6 LRB3
RB4 8 108 RB4
LRB4 108 0 LRB4
RB5 10 110 RB5
LRB5 110 0 LRB5
RB6 12 112 RB6
LRB6 112 13 LRB6
RB7 14 114 RB7
LRB7 114 15 LRB7
RB8 15 115 RB8
LRB8 115 0 LRB8
RB9 17 117 RB9
LRB9 117 0 LRB9
RB10 19 119 RB10
LRB10 119 0 LRB10
RB11 22 122 RB11
LRB11 122 15 LRB11
RB12 23 123 RB12
LRB12 123 0 LRB12
RB13 26 126 RB13
LRB13 126 0 LRB13
RB14 29 129 RB14
LRB14 129 34 LRB14
RB15 34 130 RB15
LRB15 130 31 LRB15
RB16 28 128 RB16
LRB16 128 33 LRB16
RB17 35 135 RB17
LRB17 135 0 LRB17
RB18 37 137 RB18
LRB18 137 0 LRB18
.ends LSMITLL_XNOR

*$Ports  a b clk q
.subckt LSMITLL_XNORT a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7

.param B1=2.0
.param B2=2.74
.param B3=2.23
.param B4=B1
.param B5=B2
.param B6=B3
.param B7=2.40
.param B8=3.29
.param B9=2.0
.param B10=2.42
.param B11=1.36
.param B12=2.40
.param B13=2.28
.param B14=1.75
.param B15=1.07
.param B16=1.54
.param B17=1.64
.param B18=2.5

.param IB1=195E-6
.param IB2=168E-6
.param IB3=IB1
.param IB4=IB2
.param IB5=175E-6
.param IB6=195E-6
.param IB7=60E-6
.param IB8=262E-6
.param IB9=53E-6
.param IB10=175E-6

.param L1=Lptl
.param L2=2.10e-12
.param L3=1p
.param L4=4.12e-12
.param L5=L1
.param L6=L2
.param L7=L3
.param L8=L4
.param L9=1p
.param L10=Lptl
.param L11=3.11e-12
.param L12=1.07E-12
.param L13=1.01E-12
.param L14=2.45e-12
.param L15=1.83e-12
.param L16=1.12e-12
.param L17=4.32e-12
.param L18=1.6p
.param L20=1.06E-12
.param L21=0.55E-12
.param L22=5.40e-12
.param L23=1.18e-12
.param L24=2.78e-12
.param L25=Lptl

.param RD=1.36

.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3          
.param RB4=B0Rs/B4         
.param RB5=B0Rs/B5         
.param RB6=B0Rs/B6          
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8         
.param RB9=B0Rs/B9         
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15
.param RB16=B0Rs/B16
.param RB17=B0Rs/B17
.param RB18=B0Rs/B18
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet
.param LRB13=(RB13/Rsheet)*Lsheet
.param LRB14=(RB14/Rsheet)*Lsheet
.param LRB15=(RB15/Rsheet)*Lsheet
.param LRB16=(RB16/Rsheet)*Lsheet
.param LRB17=(RB17/Rsheet)*Lsheet
.param LRB18=(RB18/Rsheet)*Lsheet

B1 1 2 jjmit area=B1
B2 3 4 jjmit area=B2
B3 5 6 jjmit area=B3
B4 8 9 jjmit area=B4
B5 10 11 jjmit area=B5
B6 12 13 jjmit area=B6
B7 14 15 jjmit area=B7
B8 15 16 jjmit area=B8
B9 17 18 jjmit area=B9
B10 19 20 jjmit area=B10
B11 22 15 jjmit area=B11
B12 23 24 jjmit area=B12
B13 26 27 jjmit area=B13
B14 29 34 jjmit area=B14
B15 34 31 jjmit area=B15
B16 28 33 jjmit area=B16
B17 35 36 jjmit area=B17
B18 37 38 jjmit area=B18

LP1 2 0 LP
LP2 4 0 LP
LP4 9 0 LP
LP5 11 0 LP
LP8 16 0 LP
LP9 18 0 LP
LP10 20 0 LP
LP12 24 0 LP
LP13 27 0 LP
LP17 36 0 LP
LP18 38 0 LP

IB1 0 1 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 8 pwl(0 0 5p IB3)
IB4 0 13 pwl(0 0 5p IB4)
IB5 0 17 pwl(0 0 5p IB5)
IB6 0 19 pwl(0 0 5p IB6)
IB7 0 25 pwl(0 0 5p IB7)
IB8 0 34 pwl(0 0 5p IB8)
IB9 0 35 pwl(0 0 5p IB9)
IB10 0 37 pwl(0 0 5p IB10)

L1 a 1 L1
L2 1 3 L2
L3 3 5 L3
L4 6 7 L4
L5 b 8 L5
L6 8 10 L6
L7 10 12 L7
L8 13 7 L8
L9 7 14 L9
L10 clk 17 L10
L11 17 19 L11
L12 19 21 L12
L13 21 22 L13
L14 21 23 L14
L15 23 25 L15
L16 25 26 L16
L17 26 28 L17
L18 15 29 L18
L20 31 32 L20
L21 33 32 L21
L22 34 28 L22
L23 32 35 L23
L24 35 37 L24
L25 37 39 L25
RD 39 q RD

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 3 103 RB2
LRB2 103 0 LRB2
RB3 5 105 RB3
LRB3 105 6 LRB3
RB4 8 108 RB4
LRB4 108 0 LRB4
RB5 10 110 RB5
LRB5 110 0 LRB5
RB6 12 112 RB6
LRB6 112 13 LRB6
RB7 14 114 RB7
LRB7 114 15 LRB7
RB8 15 115 RB8
LRB8 115 0 LRB8
RB9 17 117 RB9
LRB9 117 0 LRB9
RB10 19 119 RB10
LRB10 119 0 LRB10
RB11 22 122 RB11
LRB11 122 15 LRB11
RB12 23 123 RB12
LRB12 123 0 LRB12
RB13 26 126 RB13
LRB13 126 0 LRB13
RB14 29 129 RB14
LRB14 129 34 LRB14
RB15 34 130 RB15
LRB15 130 31 LRB15
RB16 28 128 RB16
LRB16 128 33 LRB16
RB17 35 135 RB17
LRB17 135 0 LRB17
RB18 37 137 RB18
LRB18 137 0 LRB18
.ends LSMITLL_XNORT

