.subckt 1_to_3_split a q0 q1 q2 
XSPLIT0 LSmitll_SPLIT a  a0 a1 
XSPLIT1 LSmitll_SPLIT a0 q0 q1 
XSPLIT2 LSMITLL_BUFF  a1 q2
.ends 1_to_3_split

* 1 to 4 clock splitter
.subckt 1_to_4_split a q0 q1 q2 q3
XSPLIT0 LSmitll_SPLIT a  a0 a1 
XSPLIT1 LSmitll_SPLIT a0 q0 q1 
XSPLIT2 LSmitll_SPLIT a1 q2 q3
.ends 1_to_4_split

.subckt 1_to_5_split a q0 q1 q2 q3 q4
XSPLIT0 LSmitll_SPLIT a  a0   a1 
XSPLIT1 LSmitll_SPLIT a0 a0_0 a0_1
XSPLIT2 LSmitll_SPLIT a1 a1_0 a1_1
XBUFF0 LSMITLL_BUFF a0_0 q0
XBUFF1 LSMITLL_BUFF a0_1 q1
XBUFF2 LSMITLL_BUFF a1_0 q2
XSPLIT3 LSmitll_SPLIT a1_1 q3 q4
.ends 1_to_5_split

.subckt 1_to_6_split a q0 q1 q2 q3 q4 q5
XSPLIT0 LSmitll_SPLIT a  a0   a1 
XSPLIT1 LSmitll_SPLIT a0 a0_0 a0_1
XSPLIT2 LSmitll_SPLIT a1 a1_0 a1_1
XBUFF0 LSMITLL_BUFF a0_0 q0
XBUFF1 LSMITLL_BUFF a0_1 q1
XBUFF2 LSmitll_SPLIT a1_0 q2 q3
XSPLIT3 LSmitll_SPLIT a1_1 q4 q5
.ends 1_to_6_split

* 1 to 8 clock splitter
.subckt 1_to_8_split a q0 q1 q2 q3 q4 q5 q6 q7
XSPLIT0 LSmitll_SPLIT a a0 a1 
XSPLIT1 LSmitll_SPLIT a0 a0_0 a0_1
XSPLIT2 LSmitll_SPLIT a1 a1_0 a1_1
XSPLIT3 LSmitll_SPLIT a0_0 q0 q1
XSPLIT4 LSmitll_SPLIT a0_1 q2 q3
XSPLIT5 LSmitll_SPLIT a1_0 q4 q5
XSPLIT6 LSmitll_SPLIT a1_1 q6 q7
.ends 1_to_8_split

* 1 to 16 clock splitter
.subckt 1_to_16_split a q0 q1 q2 q3 q4 q5 q6 q7 q8 q9 q10 q11 q12 q13 q14 q15
XSPLIT0  LSmitll_SPLIT a a0 a1
XSPLIT1  LSmitll_SPLIT a0 a0_0 a0_1
XSPLIT2  LSmitll_SPLIT a1 a1_0 a1_1
XSPLIT3  LSmitll_SPLIT a0_0 a0_0_0 a0_0_1
XSPLIT4  LSmitll_SPLIT a0_1 a0_1_0 a0_1_1
XSPLIT5  LSmitll_SPLIT a1_0 a1_0_0 a1_0_1
XSPLIT6  LSmitll_SPLIT a1_1 a1_1_0 a1_1_1
XSPLIT7  LSmitll_SPLIT a0_0_0 q0 q1
XSPLIT8  LSmitll_SPLIT a0_0_1 q2 q3
XSPLIT9  LSmitll_SPLIT a0_1_0 q4 q5 
XSPLIT10 LSmitll_SPLIT a0_1_1 q6 q7
XSPLIT11 LSmitll_SPLIT a1_0_0 q8 q9
XSPLIT12 LSmitll_SPLIT a1_0_1 q10 q11
XSPLIT13 LSmitll_SPLIT a1_1_0 q12 q13
XSPLIT14 LSmitll_SPLIT a1_1_1 q14 q15
.ends 1_to_16_split

* 1 to 32 clock splitter
.subckt 1_to_32_split a q0 q1 q2 q3 q4 q5 q6 q7 q8 q9 q10 q11 q12 q13 q14 q15 q16 q17 q18 q19 q20 q21 q22 q23 q24 q25 q26 q27 q28 q29 q30 q31 
XSPLIT_16 1_to_16_split a 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 
XSPLIT1 LSmitll_SPLIT 1 q0 q1
XSPLIT2 LSmitll_SPLIT 2 q2 q3
XSPLIT3 LSmitll_SPLIT 3 q4 q5
XSPLIT4 LSmitll_SPLIT 4 q6 q7
XSPLIT5 LSmitll_SPLIT 5 q8 q9
XSPLIT6 LSmitll_SPLIT 6 q10 q11
XSPLIT7 LSmitll_SPLIT 7 q12 q13
XSPLIT8 LSmitll_SPLIT 8 q14 q15
XSPLIT9 LSmitll_SPLIT 9 q16 q17
XSPLIT10 LSmitll_SPLIT 10 q18 q19
XSPLIT11 LSmitll_SPLIT 11 q20 q21
XSPLIT12 LSmitll_SPLIT 12 q22 q23
XSPLIT13 LSmitll_SPLIT 13 q24 q25
XSPLIT14 LSmitll_SPLIT 14 q26 q27
XSPLIT15 LSmitll_SPLIT 15 q28 q29
XSPLIT16 LSmitll_SPLIT 16 q30 q31
.ends 1_to_32_split

* 1 to 64 clock splitter
.subckt 1_to_64_split a q0 q1 q2 q3 q4 q5 q6 q7 q8 q9 q10 q11 q12 q13 q14 q15 q16 q17 q18 q19 q20 q21 q22 q23 q24 q25 q26 q27 q28 q29 q30 q31 q32 q33 q34 q35 q36 q37 q38 q39 q40 q41 q42 q43 q44 q45 q46 q47 q48 q49 q50 q51 q52 q53 q54 q55 q56 q57 q58 q59 q60 q61 q62 q63 
XSPLIT_32 1_to_32_split a 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 
XSPLIT1 LSmitll_SPLIT 1 q0 q1
XSPLIT2 LSmitll_SPLIT 2 q2 q3
XSPLIT3 LSmitll_SPLIT 3 q4 q5
XSPLIT4 LSmitll_SPLIT 4 q6 q7
XSPLIT5 LSmitll_SPLIT 5 q8 q9
XSPLIT6 LSmitll_SPLIT 6 q10 q11
XSPLIT7 LSmitll_SPLIT 7 q12 q13
XSPLIT8 LSmitll_SPLIT 8 q14 q15
XSPLIT9 LSmitll_SPLIT 9 q16 q17
XSPLIT10 LSmitll_SPLIT 10 q18 q19
XSPLIT11 LSmitll_SPLIT 11 q20 q21
XSPLIT12 LSmitll_SPLIT 12 q22 q23
XSPLIT13 LSmitll_SPLIT 13 q24 q25
XSPLIT14 LSmitll_SPLIT 14 q26 q27
XSPLIT15 LSmitll_SPLIT 15 q28 q29
XSPLIT16 LSmitll_SPLIT 16 q30 q31
XSPLIT17 LSmitll_SPLIT 17 q32 q33
XSPLIT18 LSmitll_SPLIT 18 q34 q35
XSPLIT19 LSmitll_SPLIT 19 q36 q37
XSPLIT20 LSmitll_SPLIT 20 q38 q39
XSPLIT21 LSmitll_SPLIT 21 q40 q41
XSPLIT22 LSmitll_SPLIT 22 q42 q43
XSPLIT23 LSmitll_SPLIT 23 q44 q45
XSPLIT24 LSmitll_SPLIT 24 q46 q47
XSPLIT25 LSmitll_SPLIT 25 q48 q49
XSPLIT26 LSmitll_SPLIT 26 q50 q51
XSPLIT27 LSmitll_SPLIT 27 q52 q53
XSPLIT28 LSmitll_SPLIT 28 q54 q55
XSPLIT29 LSmitll_SPLIT 29 q56 q57
XSPLIT30 LSmitll_SPLIT 30 q58 q59
XSPLIT31 LSmitll_SPLIT 31 q60 q61
XSPLIT32 LSmitll_SPLIT 32 q62 q63
.ends 1_to_64_split

.subckt 1_to_128_split a q0 q1 q2 q3 q4 q5 q6 q7 q8 q9 q10 q11 q12 q13 q14 q15 q16 q17 q18 q19 q20 q21 q22 q23 q24 q25 q26 q27 q28 q29 q30 q31 q32 q33 q34 q35 q36 q37 q38 q39 q40 q41 q42 q43 q44 q45 q46 q47 q48 q49 q50 q51 q52 q53 q54 q55 q56 q57 q58 q59 q60 q61 q62 q63 q64 q65 q66 q67 q68 q69 q70 q71 q72 q73 q74 q75 q76 q77 q78 q79 q80 q81 q82 q83 q84 q85 q86 q87 q88 q89 q90 q91 q92 q93 q94 q95 q96 q97 q98 q99 q100 q101 q102 q103 q104 q105 q106 q107 q108 q109 q110 q111 q112 q113 q114 q115 q116 q117 q118 q119 q120 q121 q122 q123 q124 q125 q126 q127 
XSPLIT_64 1_to_64_split a 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 
XSPLIT1 LSmitll_SPLIT 1 q0 q1
XSPLIT2 LSmitll_SPLIT 2 q2 q3
XSPLIT3 LSmitll_SPLIT 3 q4 q5
XSPLIT4 LSmitll_SPLIT 4 q6 q7
XSPLIT5 LSmitll_SPLIT 5 q8 q9
XSPLIT6 LSmitll_SPLIT 6 q10 q11
XSPLIT7 LSmitll_SPLIT 7 q12 q13
XSPLIT8 LSmitll_SPLIT 8 q14 q15
XSPLIT9 LSmitll_SPLIT 9 q16 q17
XSPLIT10 LSmitll_SPLIT 10 q18 q19
XSPLIT11 LSmitll_SPLIT 11 q20 q21
XSPLIT12 LSmitll_SPLIT 12 q22 q23
XSPLIT13 LSmitll_SPLIT 13 q24 q25
XSPLIT14 LSmitll_SPLIT 14 q26 q27
XSPLIT15 LSmitll_SPLIT 15 q28 q29
XSPLIT16 LSmitll_SPLIT 16 q30 q31
XSPLIT17 LSmitll_SPLIT 17 q32 q33
XSPLIT18 LSmitll_SPLIT 18 q34 q35
XSPLIT19 LSmitll_SPLIT 19 q36 q37
XSPLIT20 LSmitll_SPLIT 20 q38 q39
XSPLIT21 LSmitll_SPLIT 21 q40 q41
XSPLIT22 LSmitll_SPLIT 22 q42 q43
XSPLIT23 LSmitll_SPLIT 23 q44 q45
XSPLIT24 LSmitll_SPLIT 24 q46 q47
XSPLIT25 LSmitll_SPLIT 25 q48 q49
XSPLIT26 LSmitll_SPLIT 26 q50 q51
XSPLIT27 LSmitll_SPLIT 27 q52 q53
XSPLIT28 LSmitll_SPLIT 28 q54 q55
XSPLIT29 LSmitll_SPLIT 29 q56 q57
XSPLIT30 LSmitll_SPLIT 30 q58 q59
XSPLIT31 LSmitll_SPLIT 31 q60 q61
XSPLIT32 LSmitll_SPLIT 32 q62 q63
XSPLIT33 LSmitll_SPLIT 33 q64 q65
XSPLIT34 LSmitll_SPLIT 34 q66 q67
XSPLIT35 LSmitll_SPLIT 35 q68 q69
XSPLIT36 LSmitll_SPLIT 36 q70 q71
XSPLIT37 LSmitll_SPLIT 37 q72 q73
XSPLIT38 LSmitll_SPLIT 38 q74 q75
XSPLIT39 LSmitll_SPLIT 39 q76 q77
XSPLIT40 LSmitll_SPLIT 40 q78 q79
XSPLIT41 LSmitll_SPLIT 41 q80 q81
XSPLIT42 LSmitll_SPLIT 42 q82 q83
XSPLIT43 LSmitll_SPLIT 43 q84 q85
XSPLIT44 LSmitll_SPLIT 44 q86 q87
XSPLIT45 LSmitll_SPLIT 45 q88 q89
XSPLIT46 LSmitll_SPLIT 46 q90 q91
XSPLIT47 LSmitll_SPLIT 47 q92 q93
XSPLIT48 LSmitll_SPLIT 48 q94 q95
XSPLIT49 LSmitll_SPLIT 49 q96 q97
XSPLIT50 LSmitll_SPLIT 50 q98 q99
XSPLIT51 LSmitll_SPLIT 51 q100 q101
XSPLIT52 LSmitll_SPLIT 52 q102 q103
XSPLIT53 LSmitll_SPLIT 53 q104 q105
XSPLIT54 LSmitll_SPLIT 54 q106 q107
XSPLIT55 LSmitll_SPLIT 55 q108 q109
XSPLIT56 LSmitll_SPLIT 56 q110 q111
XSPLIT57 LSmitll_SPLIT 57 q112 q113
XSPLIT58 LSmitll_SPLIT 58 q114 q115
XSPLIT59 LSmitll_SPLIT 59 q116 q117
XSPLIT60 LSmitll_SPLIT 60 q118 q119
XSPLIT61 LSmitll_SPLIT 61 q120 q121
XSPLIT62 LSmitll_SPLIT 62 q122 q123
XSPLIT63 LSmitll_SPLIT 63 q124 q125
XSPLIT64 LSmitll_SPLIT 64 q126 q127
.ends 1_to_128_split

.subckt 1_to_256_split a q0 q1 q2 q3 q4 q5 q6 q7 q8 q9 q10 q11 q12 q13 q14 q15 q16 q17 q18 q19 q20 q21 q22 q23 q24 q25 q26 q27 q28 q29 q30 q31 q32 q33 q34 q35 q36 q37 q38 q39 q40 q41 q42 q43 q44 q45 q46 q47 q48 q49 q50 q51 q52 q53 q54 q55 q56 q57 q58 q59 q60 q61 q62 q63 q64 q65 q66 q67 q68 q69 q70 q71 q72 q73 q74 q75 q76 q77 q78 q79 q80 q81 q82 q83 q84 q85 q86 q87 q88 q89 q90 q91 q92 q93 q94 q95 q96 q97 q98 q99 q100 q101 q102 q103 q104 q105 q106 q107 q108 q109 q110 q111 q112 q113 q114 q115 q116 q117 q118 q119 q120 q121 q122 q123 q124 q125 q126 q127 q128 q129 q130 q131 q132 q133 q134 q135 q136 q137 q138 q139 q140 q141 q142 q143 q144 q145 q146 q147 q148 q149 q150 q151 q152 q153 q154 q155 q156 q157 q158 q159 q160 q161 q162 q163 q164 q165 q166 q167 q168 q169 q170 q171 q172 q173 q174 q175 q176 q177 q178 q179 q180 q181 q182 q183 q184 q185 q186 q187 q188 q189 q190 q191 q192 q193 q194 q195 q196 q197 q198 q199 q200 q201 q202 q203 q204 q205 q206 q207 q208 q209 q210 q211 q212 q213 q214 q215 q216 q217 q218 q219 q220 q221 q222 q223 q224 q225 q226 q227 q228 q229 q230 q231 q232 q233 q234 q235 q236 q237 q238 q239 q240 q241 q242 q243 q244 q245 q246 q247 q248 q249 q250 q251 q252 q253 q254 q255 
XSPLIT_128 1_to_128_split a 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 
XSPLIT1 LSmitll_SPLIT 1 q0 q1
XSPLIT2 LSmitll_SPLIT 2 q2 q3
XSPLIT3 LSmitll_SPLIT 3 q4 q5
XSPLIT4 LSmitll_SPLIT 4 q6 q7
XSPLIT5 LSmitll_SPLIT 5 q8 q9
XSPLIT6 LSmitll_SPLIT 6 q10 q11
XSPLIT7 LSmitll_SPLIT 7 q12 q13
XSPLIT8 LSmitll_SPLIT 8 q14 q15
XSPLIT9 LSmitll_SPLIT 9 q16 q17
XSPLIT10 LSmitll_SPLIT 10 q18 q19
XSPLIT11 LSmitll_SPLIT 11 q20 q21
XSPLIT12 LSmitll_SPLIT 12 q22 q23
XSPLIT13 LSmitll_SPLIT 13 q24 q25
XSPLIT14 LSmitll_SPLIT 14 q26 q27
XSPLIT15 LSmitll_SPLIT 15 q28 q29
XSPLIT16 LSmitll_SPLIT 16 q30 q31
XSPLIT17 LSmitll_SPLIT 17 q32 q33
XSPLIT18 LSmitll_SPLIT 18 q34 q35
XSPLIT19 LSmitll_SPLIT 19 q36 q37
XSPLIT20 LSmitll_SPLIT 20 q38 q39
XSPLIT21 LSmitll_SPLIT 21 q40 q41
XSPLIT22 LSmitll_SPLIT 22 q42 q43
XSPLIT23 LSmitll_SPLIT 23 q44 q45
XSPLIT24 LSmitll_SPLIT 24 q46 q47
XSPLIT25 LSmitll_SPLIT 25 q48 q49
XSPLIT26 LSmitll_SPLIT 26 q50 q51
XSPLIT27 LSmitll_SPLIT 27 q52 q53
XSPLIT28 LSmitll_SPLIT 28 q54 q55
XSPLIT29 LSmitll_SPLIT 29 q56 q57
XSPLIT30 LSmitll_SPLIT 30 q58 q59
XSPLIT31 LSmitll_SPLIT 31 q60 q61
XSPLIT32 LSmitll_SPLIT 32 q62 q63
XSPLIT33 LSmitll_SPLIT 33 q64 q65
XSPLIT34 LSmitll_SPLIT 34 q66 q67
XSPLIT35 LSmitll_SPLIT 35 q68 q69
XSPLIT36 LSmitll_SPLIT 36 q70 q71
XSPLIT37 LSmitll_SPLIT 37 q72 q73
XSPLIT38 LSmitll_SPLIT 38 q74 q75
XSPLIT39 LSmitll_SPLIT 39 q76 q77
XSPLIT40 LSmitll_SPLIT 40 q78 q79
XSPLIT41 LSmitll_SPLIT 41 q80 q81
XSPLIT42 LSmitll_SPLIT 42 q82 q83
XSPLIT43 LSmitll_SPLIT 43 q84 q85
XSPLIT44 LSmitll_SPLIT 44 q86 q87
XSPLIT45 LSmitll_SPLIT 45 q88 q89
XSPLIT46 LSmitll_SPLIT 46 q90 q91
XSPLIT47 LSmitll_SPLIT 47 q92 q93
XSPLIT48 LSmitll_SPLIT 48 q94 q95
XSPLIT49 LSmitll_SPLIT 49 q96 q97
XSPLIT50 LSmitll_SPLIT 50 q98 q99
XSPLIT51 LSmitll_SPLIT 51 q100 q101
XSPLIT52 LSmitll_SPLIT 52 q102 q103
XSPLIT53 LSmitll_SPLIT 53 q104 q105
XSPLIT54 LSmitll_SPLIT 54 q106 q107
XSPLIT55 LSmitll_SPLIT 55 q108 q109
XSPLIT56 LSmitll_SPLIT 56 q110 q111
XSPLIT57 LSmitll_SPLIT 57 q112 q113
XSPLIT58 LSmitll_SPLIT 58 q114 q115
XSPLIT59 LSmitll_SPLIT 59 q116 q117
XSPLIT60 LSmitll_SPLIT 60 q118 q119
XSPLIT61 LSmitll_SPLIT 61 q120 q121
XSPLIT62 LSmitll_SPLIT 62 q122 q123
XSPLIT63 LSmitll_SPLIT 63 q124 q125
XSPLIT64 LSmitll_SPLIT 64 q126 q127
XSPLIT65 LSmitll_SPLIT 65 q128 q129
XSPLIT66 LSmitll_SPLIT 66 q130 q131
XSPLIT67 LSmitll_SPLIT 67 q132 q133
XSPLIT68 LSmitll_SPLIT 68 q134 q135
XSPLIT69 LSmitll_SPLIT 69 q136 q137
XSPLIT70 LSmitll_SPLIT 70 q138 q139
XSPLIT71 LSmitll_SPLIT 71 q140 q141
XSPLIT72 LSmitll_SPLIT 72 q142 q143
XSPLIT73 LSmitll_SPLIT 73 q144 q145
XSPLIT74 LSmitll_SPLIT 74 q146 q147
XSPLIT75 LSmitll_SPLIT 75 q148 q149
XSPLIT76 LSmitll_SPLIT 76 q150 q151
XSPLIT77 LSmitll_SPLIT 77 q152 q153
XSPLIT78 LSmitll_SPLIT 78 q154 q155
XSPLIT79 LSmitll_SPLIT 79 q156 q157
XSPLIT80 LSmitll_SPLIT 80 q158 q159
XSPLIT81 LSmitll_SPLIT 81 q160 q161
XSPLIT82 LSmitll_SPLIT 82 q162 q163
XSPLIT83 LSmitll_SPLIT 83 q164 q165
XSPLIT84 LSmitll_SPLIT 84 q166 q167
XSPLIT85 LSmitll_SPLIT 85 q168 q169
XSPLIT86 LSmitll_SPLIT 86 q170 q171
XSPLIT87 LSmitll_SPLIT 87 q172 q173
XSPLIT88 LSmitll_SPLIT 88 q174 q175
XSPLIT89 LSmitll_SPLIT 89 q176 q177
XSPLIT90 LSmitll_SPLIT 90 q178 q179
XSPLIT91 LSmitll_SPLIT 91 q180 q181
XSPLIT92 LSmitll_SPLIT 92 q182 q183
XSPLIT93 LSmitll_SPLIT 93 q184 q185
XSPLIT94 LSmitll_SPLIT 94 q186 q187
XSPLIT95 LSmitll_SPLIT 95 q188 q189
XSPLIT96 LSmitll_SPLIT 96 q190 q191
XSPLIT97 LSmitll_SPLIT 97 q192 q193
XSPLIT98 LSmitll_SPLIT 98 q194 q195
XSPLIT99 LSmitll_SPLIT 99 q196 q197
XSPLIT100 LSmitll_SPLIT 100 q198 q199
XSPLIT101 LSmitll_SPLIT 101 q200 q201
XSPLIT102 LSmitll_SPLIT 102 q202 q203
XSPLIT103 LSmitll_SPLIT 103 q204 q205
XSPLIT104 LSmitll_SPLIT 104 q206 q207
XSPLIT105 LSmitll_SPLIT 105 q208 q209
XSPLIT106 LSmitll_SPLIT 106 q210 q211
XSPLIT107 LSmitll_SPLIT 107 q212 q213
XSPLIT108 LSmitll_SPLIT 108 q214 q215
XSPLIT109 LSmitll_SPLIT 109 q216 q217
XSPLIT110 LSmitll_SPLIT 110 q218 q219
XSPLIT111 LSmitll_SPLIT 111 q220 q221
XSPLIT112 LSmitll_SPLIT 112 q222 q223
XSPLIT113 LSmitll_SPLIT 113 q224 q225
XSPLIT114 LSmitll_SPLIT 114 q226 q227
XSPLIT115 LSmitll_SPLIT 115 q228 q229
XSPLIT116 LSmitll_SPLIT 116 q230 q231
XSPLIT117 LSmitll_SPLIT 117 q232 q233
XSPLIT118 LSmitll_SPLIT 118 q234 q235
XSPLIT119 LSmitll_SPLIT 119 q236 q237
XSPLIT120 LSmitll_SPLIT 120 q238 q239
XSPLIT121 LSmitll_SPLIT 121 q240 q241
XSPLIT122 LSmitll_SPLIT 122 q242 q243
XSPLIT123 LSmitll_SPLIT 123 q244 q245
XSPLIT124 LSmitll_SPLIT 124 q246 q247
XSPLIT125 LSmitll_SPLIT 125 q248 q249
XSPLIT126 LSmitll_SPLIT 126 q250 q251
XSPLIT127 LSmitll_SPLIT 127 q252 q253
XSPLIT128 LSmitll_SPLIT 128 q254 q255
.ends 1_to_256_split

.subckt 1_to_512_split a q0 q1 q2 q3 q4 q5 q6 q7 q8 q9 q10 q11 q12 q13 q14 q15 q16 q17 q18 q19 q20 q21 q22 q23 q24 q25 q26 q27 q28 q29 q30 q31 q32 q33 q34 q35 q36 q37 q38 q39 q40 q41 q42 q43 q44 q45 q46 q47 q48 q49 q50 q51 q52 q53 q54 q55 q56 q57 q58 q59 q60 q61 q62 q63 q64 q65 q66 q67 q68 q69 q70 q71 q72 q73 q74 q75 q76 q77 q78 q79 q80 q81 q82 q83 q84 q85 q86 q87 q88 q89 q90 q91 q92 q93 q94 q95 q96 q97 q98 q99 q100 q101 q102 q103 q104 q105 q106 q107 q108 q109 q110 q111 q112 q113 q114 q115 q116 q117 q118 q119 q120 q121 q122 q123 q124 q125 q126 q127 q128 q129 q130 q131 q132 q133 q134 q135 q136 q137 q138 q139 q140 q141 q142 q143 q144 q145 q146 q147 q148 q149 q150 q151 q152 q153 q154 q155 q156 q157 q158 q159 q160 q161 q162 q163 q164 q165 q166 q167 q168 q169 q170 q171 q172 q173 q174 q175 q176 q177 q178 q179 q180 q181 q182 q183 q184 q185 q186 q187 q188 q189 q190 q191 q192 q193 q194 q195 q196 q197 q198 q199 q200 q201 q202 q203 q204 q205 q206 q207 q208 q209 q210 q211 q212 q213 q214 q215 q216 q217 q218 q219 q220 q221 q222 q223 q224 q225 q226 q227 q228 q229 q230 q231 q232 q233 q234 q235 q236 q237 q238 q239 q240 q241 q242 q243 q244 q245 q246 q247 q248 q249 q250 q251 q252 q253 q254 q255 q256 q257 q258 q259 q260 q261 q262 q263 q264 q265 q266 q267 q268 q269 q270 q271 q272 q273 q274 q275 q276 q277 q278 q279 q280 q281 q282 q283 q284 q285 q286 q287 q288 q289 q290 q291 q292 q293 q294 q295 q296 q297 q298 q299 q300 q301 q302 q303 q304 q305 q306 q307 q308 q309 q310 q311 q312 q313 q314 q315 q316 q317 q318 q319 q320 q321 q322 q323 q324 q325 q326 q327 q328 q329 q330 q331 q332 q333 q334 q335 q336 q337 q338 q339 q340 q341 q342 q343 q344 q345 q346 q347 q348 q349 q350 q351 q352 q353 q354 q355 q356 q357 q358 q359 q360 q361 q362 q363 q364 q365 q366 q367 q368 q369 q370 q371 q372 q373 q374 q375 q376 q377 q378 q379 q380 q381 q382 q383 q384 q385 q386 q387 q388 q389 q390 q391 q392 q393 q394 q395 q396 q397 q398 q399 q400 q401 q402 q403 q404 q405 q406 q407 q408 q409 q410 q411 q412 q413 q414 q415 q416 q417 q418 q419 q420 q421 q422 q423 q424 q425 q426 q427 q428 q429 q430 q431 q432 q433 q434 q435 q436 q437 q438 q439 q440 q441 q442 q443 q444 q445 q446 q447 q448 q449 q450 q451 q452 q453 q454 q455 q456 q457 q458 q459 q460 q461 q462 q463 q464 q465 q466 q467 q468 q469 q470 q471 q472 q473 q474 q475 q476 q477 q478 q479 q480 q481 q482 q483 q484 q485 q486 q487 q488 q489 q490 q491 q492 q493 q494 q495 q496 q497 q498 q499 q500 q501 q502 q503 q504 q505 q506 q507 q508 q509 q510 q511 
XSPLIT_256 1_to_256_split a 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 
XSPLIT1 LSmitll_SPLIT 1 q0 q1
XSPLIT2 LSmitll_SPLIT 2 q2 q3
XSPLIT3 LSmitll_SPLIT 3 q4 q5
XSPLIT4 LSmitll_SPLIT 4 q6 q7
XSPLIT5 LSmitll_SPLIT 5 q8 q9
XSPLIT6 LSmitll_SPLIT 6 q10 q11
XSPLIT7 LSmitll_SPLIT 7 q12 q13
XSPLIT8 LSmitll_SPLIT 8 q14 q15
XSPLIT9 LSmitll_SPLIT 9 q16 q17
XSPLIT10 LSmitll_SPLIT 10 q18 q19
XSPLIT11 LSmitll_SPLIT 11 q20 q21
XSPLIT12 LSmitll_SPLIT 12 q22 q23
XSPLIT13 LSmitll_SPLIT 13 q24 q25
XSPLIT14 LSmitll_SPLIT 14 q26 q27
XSPLIT15 LSmitll_SPLIT 15 q28 q29
XSPLIT16 LSmitll_SPLIT 16 q30 q31
XSPLIT17 LSmitll_SPLIT 17 q32 q33
XSPLIT18 LSmitll_SPLIT 18 q34 q35
XSPLIT19 LSmitll_SPLIT 19 q36 q37
XSPLIT20 LSmitll_SPLIT 20 q38 q39
XSPLIT21 LSmitll_SPLIT 21 q40 q41
XSPLIT22 LSmitll_SPLIT 22 q42 q43
XSPLIT23 LSmitll_SPLIT 23 q44 q45
XSPLIT24 LSmitll_SPLIT 24 q46 q47
XSPLIT25 LSmitll_SPLIT 25 q48 q49
XSPLIT26 LSmitll_SPLIT 26 q50 q51
XSPLIT27 LSmitll_SPLIT 27 q52 q53
XSPLIT28 LSmitll_SPLIT 28 q54 q55
XSPLIT29 LSmitll_SPLIT 29 q56 q57
XSPLIT30 LSmitll_SPLIT 30 q58 q59
XSPLIT31 LSmitll_SPLIT 31 q60 q61
XSPLIT32 LSmitll_SPLIT 32 q62 q63
XSPLIT33 LSmitll_SPLIT 33 q64 q65
XSPLIT34 LSmitll_SPLIT 34 q66 q67
XSPLIT35 LSmitll_SPLIT 35 q68 q69
XSPLIT36 LSmitll_SPLIT 36 q70 q71
XSPLIT37 LSmitll_SPLIT 37 q72 q73
XSPLIT38 LSmitll_SPLIT 38 q74 q75
XSPLIT39 LSmitll_SPLIT 39 q76 q77
XSPLIT40 LSmitll_SPLIT 40 q78 q79
XSPLIT41 LSmitll_SPLIT 41 q80 q81
XSPLIT42 LSmitll_SPLIT 42 q82 q83
XSPLIT43 LSmitll_SPLIT 43 q84 q85
XSPLIT44 LSmitll_SPLIT 44 q86 q87
XSPLIT45 LSmitll_SPLIT 45 q88 q89
XSPLIT46 LSmitll_SPLIT 46 q90 q91
XSPLIT47 LSmitll_SPLIT 47 q92 q93
XSPLIT48 LSmitll_SPLIT 48 q94 q95
XSPLIT49 LSmitll_SPLIT 49 q96 q97
XSPLIT50 LSmitll_SPLIT 50 q98 q99
XSPLIT51 LSmitll_SPLIT 51 q100 q101
XSPLIT52 LSmitll_SPLIT 52 q102 q103
XSPLIT53 LSmitll_SPLIT 53 q104 q105
XSPLIT54 LSmitll_SPLIT 54 q106 q107
XSPLIT55 LSmitll_SPLIT 55 q108 q109
XSPLIT56 LSmitll_SPLIT 56 q110 q111
XSPLIT57 LSmitll_SPLIT 57 q112 q113
XSPLIT58 LSmitll_SPLIT 58 q114 q115
XSPLIT59 LSmitll_SPLIT 59 q116 q117
XSPLIT60 LSmitll_SPLIT 60 q118 q119
XSPLIT61 LSmitll_SPLIT 61 q120 q121
XSPLIT62 LSmitll_SPLIT 62 q122 q123
XSPLIT63 LSmitll_SPLIT 63 q124 q125
XSPLIT64 LSmitll_SPLIT 64 q126 q127
XSPLIT65 LSmitll_SPLIT 65 q128 q129
XSPLIT66 LSmitll_SPLIT 66 q130 q131
XSPLIT67 LSmitll_SPLIT 67 q132 q133
XSPLIT68 LSmitll_SPLIT 68 q134 q135
XSPLIT69 LSmitll_SPLIT 69 q136 q137
XSPLIT70 LSmitll_SPLIT 70 q138 q139
XSPLIT71 LSmitll_SPLIT 71 q140 q141
XSPLIT72 LSmitll_SPLIT 72 q142 q143
XSPLIT73 LSmitll_SPLIT 73 q144 q145
XSPLIT74 LSmitll_SPLIT 74 q146 q147
XSPLIT75 LSmitll_SPLIT 75 q148 q149
XSPLIT76 LSmitll_SPLIT 76 q150 q151
XSPLIT77 LSmitll_SPLIT 77 q152 q153
XSPLIT78 LSmitll_SPLIT 78 q154 q155
XSPLIT79 LSmitll_SPLIT 79 q156 q157
XSPLIT80 LSmitll_SPLIT 80 q158 q159
XSPLIT81 LSmitll_SPLIT 81 q160 q161
XSPLIT82 LSmitll_SPLIT 82 q162 q163
XSPLIT83 LSmitll_SPLIT 83 q164 q165
XSPLIT84 LSmitll_SPLIT 84 q166 q167
XSPLIT85 LSmitll_SPLIT 85 q168 q169
XSPLIT86 LSmitll_SPLIT 86 q170 q171
XSPLIT87 LSmitll_SPLIT 87 q172 q173
XSPLIT88 LSmitll_SPLIT 88 q174 q175
XSPLIT89 LSmitll_SPLIT 89 q176 q177
XSPLIT90 LSmitll_SPLIT 90 q178 q179
XSPLIT91 LSmitll_SPLIT 91 q180 q181
XSPLIT92 LSmitll_SPLIT 92 q182 q183
XSPLIT93 LSmitll_SPLIT 93 q184 q185
XSPLIT94 LSmitll_SPLIT 94 q186 q187
XSPLIT95 LSmitll_SPLIT 95 q188 q189
XSPLIT96 LSmitll_SPLIT 96 q190 q191
XSPLIT97 LSmitll_SPLIT 97 q192 q193
XSPLIT98 LSmitll_SPLIT 98 q194 q195
XSPLIT99 LSmitll_SPLIT 99 q196 q197
XSPLIT100 LSmitll_SPLIT 100 q198 q199
XSPLIT101 LSmitll_SPLIT 101 q200 q201
XSPLIT102 LSmitll_SPLIT 102 q202 q203
XSPLIT103 LSmitll_SPLIT 103 q204 q205
XSPLIT104 LSmitll_SPLIT 104 q206 q207
XSPLIT105 LSmitll_SPLIT 105 q208 q209
XSPLIT106 LSmitll_SPLIT 106 q210 q211
XSPLIT107 LSmitll_SPLIT 107 q212 q213
XSPLIT108 LSmitll_SPLIT 108 q214 q215
XSPLIT109 LSmitll_SPLIT 109 q216 q217
XSPLIT110 LSmitll_SPLIT 110 q218 q219
XSPLIT111 LSmitll_SPLIT 111 q220 q221
XSPLIT112 LSmitll_SPLIT 112 q222 q223
XSPLIT113 LSmitll_SPLIT 113 q224 q225
XSPLIT114 LSmitll_SPLIT 114 q226 q227
XSPLIT115 LSmitll_SPLIT 115 q228 q229
XSPLIT116 LSmitll_SPLIT 116 q230 q231
XSPLIT117 LSmitll_SPLIT 117 q232 q233
XSPLIT118 LSmitll_SPLIT 118 q234 q235
XSPLIT119 LSmitll_SPLIT 119 q236 q237
XSPLIT120 LSmitll_SPLIT 120 q238 q239
XSPLIT121 LSmitll_SPLIT 121 q240 q241
XSPLIT122 LSmitll_SPLIT 122 q242 q243
XSPLIT123 LSmitll_SPLIT 123 q244 q245
XSPLIT124 LSmitll_SPLIT 124 q246 q247
XSPLIT125 LSmitll_SPLIT 125 q248 q249
XSPLIT126 LSmitll_SPLIT 126 q250 q251
XSPLIT127 LSmitll_SPLIT 127 q252 q253
XSPLIT128 LSmitll_SPLIT 128 q254 q255
XSPLIT129 LSmitll_SPLIT 129 q256 q257
XSPLIT130 LSmitll_SPLIT 130 q258 q259
XSPLIT131 LSmitll_SPLIT 131 q260 q261
XSPLIT132 LSmitll_SPLIT 132 q262 q263
XSPLIT133 LSmitll_SPLIT 133 q264 q265
XSPLIT134 LSmitll_SPLIT 134 q266 q267
XSPLIT135 LSmitll_SPLIT 135 q268 q269
XSPLIT136 LSmitll_SPLIT 136 q270 q271
XSPLIT137 LSmitll_SPLIT 137 q272 q273
XSPLIT138 LSmitll_SPLIT 138 q274 q275
XSPLIT139 LSmitll_SPLIT 139 q276 q277
XSPLIT140 LSmitll_SPLIT 140 q278 q279
XSPLIT141 LSmitll_SPLIT 141 q280 q281
XSPLIT142 LSmitll_SPLIT 142 q282 q283
XSPLIT143 LSmitll_SPLIT 143 q284 q285
XSPLIT144 LSmitll_SPLIT 144 q286 q287
XSPLIT145 LSmitll_SPLIT 145 q288 q289
XSPLIT146 LSmitll_SPLIT 146 q290 q291
XSPLIT147 LSmitll_SPLIT 147 q292 q293
XSPLIT148 LSmitll_SPLIT 148 q294 q295
XSPLIT149 LSmitll_SPLIT 149 q296 q297
XSPLIT150 LSmitll_SPLIT 150 q298 q299
XSPLIT151 LSmitll_SPLIT 151 q300 q301
XSPLIT152 LSmitll_SPLIT 152 q302 q303
XSPLIT153 LSmitll_SPLIT 153 q304 q305
XSPLIT154 LSmitll_SPLIT 154 q306 q307
XSPLIT155 LSmitll_SPLIT 155 q308 q309
XSPLIT156 LSmitll_SPLIT 156 q310 q311
XSPLIT157 LSmitll_SPLIT 157 q312 q313
XSPLIT158 LSmitll_SPLIT 158 q314 q315
XSPLIT159 LSmitll_SPLIT 159 q316 q317
XSPLIT160 LSmitll_SPLIT 160 q318 q319
XSPLIT161 LSmitll_SPLIT 161 q320 q321
XSPLIT162 LSmitll_SPLIT 162 q322 q323
XSPLIT163 LSmitll_SPLIT 163 q324 q325
XSPLIT164 LSmitll_SPLIT 164 q326 q327
XSPLIT165 LSmitll_SPLIT 165 q328 q329
XSPLIT166 LSmitll_SPLIT 166 q330 q331
XSPLIT167 LSmitll_SPLIT 167 q332 q333
XSPLIT168 LSmitll_SPLIT 168 q334 q335
XSPLIT169 LSmitll_SPLIT 169 q336 q337
XSPLIT170 LSmitll_SPLIT 170 q338 q339
XSPLIT171 LSmitll_SPLIT 171 q340 q341
XSPLIT172 LSmitll_SPLIT 172 q342 q343
XSPLIT173 LSmitll_SPLIT 173 q344 q345
XSPLIT174 LSmitll_SPLIT 174 q346 q347
XSPLIT175 LSmitll_SPLIT 175 q348 q349
XSPLIT176 LSmitll_SPLIT 176 q350 q351
XSPLIT177 LSmitll_SPLIT 177 q352 q353
XSPLIT178 LSmitll_SPLIT 178 q354 q355
XSPLIT179 LSmitll_SPLIT 179 q356 q357
XSPLIT180 LSmitll_SPLIT 180 q358 q359
XSPLIT181 LSmitll_SPLIT 181 q360 q361
XSPLIT182 LSmitll_SPLIT 182 q362 q363
XSPLIT183 LSmitll_SPLIT 183 q364 q365
XSPLIT184 LSmitll_SPLIT 184 q366 q367
XSPLIT185 LSmitll_SPLIT 185 q368 q369
XSPLIT186 LSmitll_SPLIT 186 q370 q371
XSPLIT187 LSmitll_SPLIT 187 q372 q373
XSPLIT188 LSmitll_SPLIT 188 q374 q375
XSPLIT189 LSmitll_SPLIT 189 q376 q377
XSPLIT190 LSmitll_SPLIT 190 q378 q379
XSPLIT191 LSmitll_SPLIT 191 q380 q381
XSPLIT192 LSmitll_SPLIT 192 q382 q383
XSPLIT193 LSmitll_SPLIT 193 q384 q385
XSPLIT194 LSmitll_SPLIT 194 q386 q387
XSPLIT195 LSmitll_SPLIT 195 q388 q389
XSPLIT196 LSmitll_SPLIT 196 q390 q391
XSPLIT197 LSmitll_SPLIT 197 q392 q393
XSPLIT198 LSmitll_SPLIT 198 q394 q395
XSPLIT199 LSmitll_SPLIT 199 q396 q397
XSPLIT200 LSmitll_SPLIT 200 q398 q399
XSPLIT201 LSmitll_SPLIT 201 q400 q401
XSPLIT202 LSmitll_SPLIT 202 q402 q403
XSPLIT203 LSmitll_SPLIT 203 q404 q405
XSPLIT204 LSmitll_SPLIT 204 q406 q407
XSPLIT205 LSmitll_SPLIT 205 q408 q409
XSPLIT206 LSmitll_SPLIT 206 q410 q411
XSPLIT207 LSmitll_SPLIT 207 q412 q413
XSPLIT208 LSmitll_SPLIT 208 q414 q415
XSPLIT209 LSmitll_SPLIT 209 q416 q417
XSPLIT210 LSmitll_SPLIT 210 q418 q419
XSPLIT211 LSmitll_SPLIT 211 q420 q421
XSPLIT212 LSmitll_SPLIT 212 q422 q423
XSPLIT213 LSmitll_SPLIT 213 q424 q425
XSPLIT214 LSmitll_SPLIT 214 q426 q427
XSPLIT215 LSmitll_SPLIT 215 q428 q429
XSPLIT216 LSmitll_SPLIT 216 q430 q431
XSPLIT217 LSmitll_SPLIT 217 q432 q433
XSPLIT218 LSmitll_SPLIT 218 q434 q435
XSPLIT219 LSmitll_SPLIT 219 q436 q437
XSPLIT220 LSmitll_SPLIT 220 q438 q439
XSPLIT221 LSmitll_SPLIT 221 q440 q441
XSPLIT222 LSmitll_SPLIT 222 q442 q443
XSPLIT223 LSmitll_SPLIT 223 q444 q445
XSPLIT224 LSmitll_SPLIT 224 q446 q447
XSPLIT225 LSmitll_SPLIT 225 q448 q449
XSPLIT226 LSmitll_SPLIT 226 q450 q451
XSPLIT227 LSmitll_SPLIT 227 q452 q453
XSPLIT228 LSmitll_SPLIT 228 q454 q455
XSPLIT229 LSmitll_SPLIT 229 q456 q457
XSPLIT230 LSmitll_SPLIT 230 q458 q459
XSPLIT231 LSmitll_SPLIT 231 q460 q461
XSPLIT232 LSmitll_SPLIT 232 q462 q463
XSPLIT233 LSmitll_SPLIT 233 q464 q465
XSPLIT234 LSmitll_SPLIT 234 q466 q467
XSPLIT235 LSmitll_SPLIT 235 q468 q469
XSPLIT236 LSmitll_SPLIT 236 q470 q471
XSPLIT237 LSmitll_SPLIT 237 q472 q473
XSPLIT238 LSmitll_SPLIT 238 q474 q475
XSPLIT239 LSmitll_SPLIT 239 q476 q477
XSPLIT240 LSmitll_SPLIT 240 q478 q479
XSPLIT241 LSmitll_SPLIT 241 q480 q481
XSPLIT242 LSmitll_SPLIT 242 q482 q483
XSPLIT243 LSmitll_SPLIT 243 q484 q485
XSPLIT244 LSmitll_SPLIT 244 q486 q487
XSPLIT245 LSmitll_SPLIT 245 q488 q489
XSPLIT246 LSmitll_SPLIT 246 q490 q491
XSPLIT247 LSmitll_SPLIT 247 q492 q493
XSPLIT248 LSmitll_SPLIT 248 q494 q495
XSPLIT249 LSmitll_SPLIT 249 q496 q497
XSPLIT250 LSmitll_SPLIT 250 q498 q499
XSPLIT251 LSmitll_SPLIT 251 q500 q501
XSPLIT252 LSmitll_SPLIT 252 q502 q503
XSPLIT253 LSmitll_SPLIT 253 q504 q505
XSPLIT254 LSmitll_SPLIT 254 q506 q507
XSPLIT255 LSmitll_SPLIT 255 q508 q509
XSPLIT256 LSmitll_SPLIT 256 q510 q511
.ends 1_to_512_split

.subckt 1_to_848_split a q0 q1 q2 q3 q4 q5 q6 q7 q8 q9 q10 q11 q12 q13 q14 q15 q16 q17 q18 q19 q20 q21 q22 q23 q24 q25 q26 q27 q28 q29 q30 q31 q32 q33 q34 q35 q36 q37 q38 q39 q40 q41 q42 q43 q44 q45 q46 q47 q48 q49 q50 q51 q52 q53 q54 q55 q56 q57 q58 q59 q60 q61 q62 q63 q64 q65 q66 q67 q68 q69 q70 q71 q72 q73 q74 q75 q76 q77 q78 q79 q80 q81 q82 q83 q84 q85 q86 q87 q88 q89 q90 q91 q92 q93 q94 q95 q96 q97 q98 q99 q100 q101 q102 q103 q104 q105 q106 q107 q108 q109 q110 q111 q112 q113 q114 q115 q116 q117 q118 q119 q120 q121 q122 q123 q124 q125 q126 q127 q128 q129 q130 q131 q132 q133 q134 q135 q136 q137 q138 q139 q140 q141 q142 q143 q144 q145 q146 q147 q148 q149 q150 q151 q152 q153 q154 q155 q156 q157 q158 q159 q160 q161 q162 q163 q164 q165 q166 q167 q168 q169 q170 q171 q172 q173 q174 q175 q176 q177 q178 q179 q180 q181 q182 q183 q184 q185 q186 q187 q188 q189 q190 q191 q192 q193 q194 q195 q196 q197 q198 q199 q200 q201 q202 q203 q204 q205 q206 q207 q208 q209 q210 q211 q212 q213 q214 q215 q216 q217 q218 q219 q220 q221 q222 q223 q224 q225 q226 q227 q228 q229 q230 q231 q232 q233 q234 q235 q236 q237 q238 q239 q240 q241 q242 q243 q244 q245 q246 q247 q248 q249 q250 q251 q252 q253 q254 q255 q256 q257 q258 q259 q260 q261 q262 q263 q264 q265 q266 q267 q268 q269 q270 q271 q272 q273 q274 q275 q276 q277 q278 q279 q280 q281 q282 q283 q284 q285 q286 q287 q288 q289 q290 q291 q292 q293 q294 q295 q296 q297 q298 q299 q300 q301 q302 q303 q304 q305 q306 q307 q308 q309 q310 q311 q312 q313 q314 q315 q316 q317 q318 q319 q320 q321 q322 q323 q324 q325 q326 q327 q328 q329 q330 q331 q332 q333 q334 q335 q336 q337 q338 q339 q340 q341 q342 q343 q344 q345 q346 q347 q348 q349 q350 q351 q352 q353 q354 q355 q356 q357 q358 q359 q360 q361 q362 q363 q364 q365 q366 q367 q368 q369 q370 q371 q372 q373 q374 q375 q376 q377 q378 q379 q380 q381 q382 q383 q384 q385 q386 q387 q388 q389 q390 q391 q392 q393 q394 q395 q396 q397 q398 q399 q400 q401 q402 q403 q404 q405 q406 q407 q408 q409 q410 q411 q412 q413 q414 q415 q416 q417 q418 q419 q420 q421 q422 q423 q424 q425 q426 q427 q428 q429 q430 q431 q432 q433 q434 q435 q436 q437 q438 q439 q440 q441 q442 q443 q444 q445 q446 q447 q448 q449 q450 q451 q452 q453 q454 q455 q456 q457 q458 q459 q460 q461 q462 q463 q464 q465 q466 q467 q468 q469 q470 q471 q472 q473 q474 q475 q476 q477 q478 q479 q480 q481 q482 q483 q484 q485 q486 q487 q488 q489 q490 q491 q492 q493 q494 q495 q496 q497 q498 q499 q500 q501 q502 q503 q504 q505 q506 q507 q508 q509 q510 q511 q512 q513 q514 q515 q516 q517 q518 q519 q520 q521 q522 q523 q524 q525 q526 q527 q528 q529 q530 q531 q532 q533 q534 q535 q536 q537 q538 q539 q540 q541 q542 q543 q544 q545 q546 q547 q548 q549 q550 q551 q552 q553 q554 q555 q556 q557 q558 q559 q560 q561 q562 q563 q564 q565 q566 q567 q568 q569 q570 q571 q572 q573 q574 q575 q576 q577 q578 q579 q580 q581 q582 q583 q584 q585 q586 q587 q588 q589 q590 q591 q592 q593 q594 q595 q596 q597 q598 q599 q600 q601 q602 q603 q604 q605 q606 q607 q608 q609 q610 q611 q612 q613 q614 q615 q616 q617 q618 q619 q620 q621 q622 q623 q624 q625 q626 q627 q628 q629 q630 q631 q632 q633 q634 q635 q636 q637 q638 q639 q640 q641 q642 q643 q644 q645 q646 q647 q648 q649 q650 q651 q652 q653 q654 q655 q656 q657 q658 q659 q660 q661 q662 q663 q664 q665 q666 q667 q668 q669 q670 q671 q672 q673 q674 q675 q676 q677 q678 q679 q680 q681 q682 q683 q684 q685 q686 q687 q688 q689 q690 q691 q692 q693 q694 q695 q696 q697 q698 q699 q700 q701 q702 q703 q704 q705 q706 q707 q708 q709 q710 q711 q712 q713 q714 q715 q716 q717 q718 q719 q720 q721 q722 q723 q724 q725 q726 q727 q728 q729 q730 q731 q732 q733 q734 q735 q736 q737 q738 q739 q740 q741 q742 q743 q744 q745 q746 q747 q748 q749 q750 q751 q752 q753 q754 q755 q756 q757 q758 q759 q760 q761 q762 q763 q764 q765 q766 q767 q768 q769 q770 q771 q772 q773 q774 q775 q776 q777 q778 q779 q780 q781 q782 q783 q784 q785 q786 q787 q788 q789 q790 q791 q792 q793 q794 q795 q796 q797 q798 q799 q800 q801 q802 q803 q804 q805 q806 q807 q808 q809 q810 q811 q812 q813 q814 q815 q816 q817 q818 q819 q820 q821 q822 q823 q824 q825 q826 q827 q828 q829 q830 q831 q832 q833 q834 q835 q836 q837 q838 q839 q840 q841 q842 q843 q844 q845 q846 q847
XSPLIT_512 1_to_512_split a 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510 511 512 
XSPLIT1 LSmitll_SPLIT 1 q0 q1
XSPLIT2 LSmitll_SPLIT 2 q2 q3
XSPLIT3 LSmitll_SPLIT 3 q4 q5
XSPLIT4 LSmitll_SPLIT 4 q6 q7
XSPLIT5 LSmitll_SPLIT 5 q8 q9
XSPLIT6 LSmitll_SPLIT 6 q10 q11
XSPLIT7 LSmitll_SPLIT 7 q12 q13
XSPLIT8 LSmitll_SPLIT 8 q14 q15
XSPLIT9 LSmitll_SPLIT 9 q16 q17
XSPLIT10 LSmitll_SPLIT 10 q18 q19
XSPLIT11 LSmitll_SPLIT 11 q20 q21
XSPLIT12 LSmitll_SPLIT 12 q22 q23
XSPLIT13 LSmitll_SPLIT 13 q24 q25
XSPLIT14 LSmitll_SPLIT 14 q26 q27
XSPLIT15 LSmitll_SPLIT 15 q28 q29
XSPLIT16 LSmitll_SPLIT 16 q30 q31
XSPLIT17 LSmitll_SPLIT 17 q32 q33
XSPLIT18 LSmitll_SPLIT 18 q34 q35
XSPLIT19 LSmitll_SPLIT 19 q36 q37
XSPLIT20 LSmitll_SPLIT 20 q38 q39
XSPLIT21 LSmitll_SPLIT 21 q40 q41
XSPLIT22 LSmitll_SPLIT 22 q42 q43
XSPLIT23 LSmitll_SPLIT 23 q44 q45
XSPLIT24 LSmitll_SPLIT 24 q46 q47
XSPLIT25 LSmitll_SPLIT 25 q48 q49
XSPLIT26 LSmitll_SPLIT 26 q50 q51
XSPLIT27 LSmitll_SPLIT 27 q52 q53
XSPLIT28 LSmitll_SPLIT 28 q54 q55
XSPLIT29 LSmitll_SPLIT 29 q56 q57
XSPLIT30 LSmitll_SPLIT 30 q58 q59
XSPLIT31 LSmitll_SPLIT 31 q60 q61
XSPLIT32 LSmitll_SPLIT 32 q62 q63
XSPLIT33 LSmitll_SPLIT 33 q64 q65
XSPLIT34 LSmitll_SPLIT 34 q66 q67
XSPLIT35 LSmitll_SPLIT 35 q68 q69
XSPLIT36 LSmitll_SPLIT 36 q70 q71
XSPLIT37 LSmitll_SPLIT 37 q72 q73
XSPLIT38 LSmitll_SPLIT 38 q74 q75
XSPLIT39 LSmitll_SPLIT 39 q76 q77
XSPLIT40 LSmitll_SPLIT 40 q78 q79
XSPLIT41 LSmitll_SPLIT 41 q80 q81
XSPLIT42 LSmitll_SPLIT 42 q82 q83
XSPLIT43 LSmitll_SPLIT 43 q84 q85
XSPLIT44 LSmitll_SPLIT 44 q86 q87
XSPLIT45 LSmitll_SPLIT 45 q88 q89
XSPLIT46 LSmitll_SPLIT 46 q90 q91
XSPLIT47 LSmitll_SPLIT 47 q92 q93
XSPLIT48 LSmitll_SPLIT 48 q94 q95
XSPLIT49 LSmitll_SPLIT 49 q96 q97
XSPLIT50 LSmitll_SPLIT 50 q98 q99
XSPLIT51 LSmitll_SPLIT 51 q100 q101
XSPLIT52 LSmitll_SPLIT 52 q102 q103
XSPLIT53 LSmitll_SPLIT 53 q104 q105
XSPLIT54 LSmitll_SPLIT 54 q106 q107
XSPLIT55 LSmitll_SPLIT 55 q108 q109
XSPLIT56 LSmitll_SPLIT 56 q110 q111
XSPLIT57 LSmitll_SPLIT 57 q112 q113
XSPLIT58 LSmitll_SPLIT 58 q114 q115
XSPLIT59 LSmitll_SPLIT 59 q116 q117
XSPLIT60 LSmitll_SPLIT 60 q118 q119
XSPLIT61 LSmitll_SPLIT 61 q120 q121
XSPLIT62 LSmitll_SPLIT 62 q122 q123
XSPLIT63 LSmitll_SPLIT 63 q124 q125
XSPLIT64 LSmitll_SPLIT 64 q126 q127
XSPLIT65 LSmitll_SPLIT 65 q128 q129
XSPLIT66 LSmitll_SPLIT 66 q130 q131
XSPLIT67 LSmitll_SPLIT 67 q132 q133
XSPLIT68 LSmitll_SPLIT 68 q134 q135
XSPLIT69 LSmitll_SPLIT 69 q136 q137
XSPLIT70 LSmitll_SPLIT 70 q138 q139
XSPLIT71 LSmitll_SPLIT 71 q140 q141
XSPLIT72 LSmitll_SPLIT 72 q142 q143
XSPLIT73 LSmitll_SPLIT 73 q144 q145
XSPLIT74 LSmitll_SPLIT 74 q146 q147
XSPLIT75 LSmitll_SPLIT 75 q148 q149
XSPLIT76 LSmitll_SPLIT 76 q150 q151
XSPLIT77 LSmitll_SPLIT 77 q152 q153
XSPLIT78 LSmitll_SPLIT 78 q154 q155
XSPLIT79 LSmitll_SPLIT 79 q156 q157
XSPLIT80 LSmitll_SPLIT 80 q158 q159
XSPLIT81 LSmitll_SPLIT 81 q160 q161
XSPLIT82 LSmitll_SPLIT 82 q162 q163
XSPLIT83 LSmitll_SPLIT 83 q164 q165
XSPLIT84 LSmitll_SPLIT 84 q166 q167
XSPLIT85 LSmitll_SPLIT 85 q168 q169
XSPLIT86 LSmitll_SPLIT 86 q170 q171
XSPLIT87 LSmitll_SPLIT 87 q172 q173
XSPLIT88 LSmitll_SPLIT 88 q174 q175
XSPLIT89 LSmitll_SPLIT 89 q176 q177
XSPLIT90 LSmitll_SPLIT 90 q178 q179
XSPLIT91 LSmitll_SPLIT 91 q180 q181
XSPLIT92 LSmitll_SPLIT 92 q182 q183
XSPLIT93 LSmitll_SPLIT 93 q184 q185
XSPLIT94 LSmitll_SPLIT 94 q186 q187
XSPLIT95 LSmitll_SPLIT 95 q188 q189
XSPLIT96 LSmitll_SPLIT 96 q190 q191
XSPLIT97 LSmitll_SPLIT 97 q192 q193
XSPLIT98 LSmitll_SPLIT 98 q194 q195
XSPLIT99 LSmitll_SPLIT 99 q196 q197
XSPLIT100 LSmitll_SPLIT 100 q198 q199
XSPLIT101 LSmitll_SPLIT 101 q200 q201
XSPLIT102 LSmitll_SPLIT 102 q202 q203
XSPLIT103 LSmitll_SPLIT 103 q204 q205
XSPLIT104 LSmitll_SPLIT 104 q206 q207
XSPLIT105 LSmitll_SPLIT 105 q208 q209
XSPLIT106 LSmitll_SPLIT 106 q210 q211
XSPLIT107 LSmitll_SPLIT 107 q212 q213
XSPLIT108 LSmitll_SPLIT 108 q214 q215
XSPLIT109 LSmitll_SPLIT 109 q216 q217
XSPLIT110 LSmitll_SPLIT 110 q218 q219
XSPLIT111 LSmitll_SPLIT 111 q220 q221
XSPLIT112 LSmitll_SPLIT 112 q222 q223
XSPLIT113 LSmitll_SPLIT 113 q224 q225
XSPLIT114 LSmitll_SPLIT 114 q226 q227
XSPLIT115 LSmitll_SPLIT 115 q228 q229
XSPLIT116 LSmitll_SPLIT 116 q230 q231
XSPLIT117 LSmitll_SPLIT 117 q232 q233
XSPLIT118 LSmitll_SPLIT 118 q234 q235
XSPLIT119 LSmitll_SPLIT 119 q236 q237
XSPLIT120 LSmitll_SPLIT 120 q238 q239
XSPLIT121 LSmitll_SPLIT 121 q240 q241
XSPLIT122 LSmitll_SPLIT 122 q242 q243
XSPLIT123 LSmitll_SPLIT 123 q244 q245
XSPLIT124 LSmitll_SPLIT 124 q246 q247
XSPLIT125 LSmitll_SPLIT 125 q248 q249
XSPLIT126 LSmitll_SPLIT 126 q250 q251
XSPLIT127 LSmitll_SPLIT 127 q252 q253
XSPLIT128 LSmitll_SPLIT 128 q254 q255
XSPLIT129 LSmitll_SPLIT 129 q256 q257
XSPLIT130 LSmitll_SPLIT 130 q258 q259
XSPLIT131 LSmitll_SPLIT 131 q260 q261
XSPLIT132 LSmitll_SPLIT 132 q262 q263
XSPLIT133 LSmitll_SPLIT 133 q264 q265
XSPLIT134 LSmitll_SPLIT 134 q266 q267
XSPLIT135 LSmitll_SPLIT 135 q268 q269
XSPLIT136 LSmitll_SPLIT 136 q270 q271
XSPLIT137 LSmitll_SPLIT 137 q272 q273
XSPLIT138 LSmitll_SPLIT 138 q274 q275
XSPLIT139 LSmitll_SPLIT 139 q276 q277
XSPLIT140 LSmitll_SPLIT 140 q278 q279
XSPLIT141 LSmitll_SPLIT 141 q280 q281
XSPLIT142 LSmitll_SPLIT 142 q282 q283
XSPLIT143 LSmitll_SPLIT 143 q284 q285
XSPLIT144 LSmitll_SPLIT 144 q286 q287
XSPLIT145 LSmitll_SPLIT 145 q288 q289
XSPLIT146 LSmitll_SPLIT 146 q290 q291
XSPLIT147 LSmitll_SPLIT 147 q292 q293
XSPLIT148 LSmitll_SPLIT 148 q294 q295
XSPLIT149 LSmitll_SPLIT 149 q296 q297
XSPLIT150 LSmitll_SPLIT 150 q298 q299
XSPLIT151 LSmitll_SPLIT 151 q300 q301
XSPLIT152 LSmitll_SPLIT 152 q302 q303
XSPLIT153 LSmitll_SPLIT 153 q304 q305
XSPLIT154 LSmitll_SPLIT 154 q306 q307
XSPLIT155 LSmitll_SPLIT 155 q308 q309
XSPLIT156 LSmitll_SPLIT 156 q310 q311
XSPLIT157 LSmitll_SPLIT 157 q312 q313
XSPLIT158 LSmitll_SPLIT 158 q314 q315
XSPLIT159 LSmitll_SPLIT 159 q316 q317
XSPLIT160 LSmitll_SPLIT 160 q318 q319
XSPLIT161 LSmitll_SPLIT 161 q320 q321
XSPLIT162 LSmitll_SPLIT 162 q322 q323
XSPLIT163 LSmitll_SPLIT 163 q324 q325
XSPLIT164 LSmitll_SPLIT 164 q326 q327
XSPLIT165 LSmitll_SPLIT 165 q328 q329
XSPLIT166 LSmitll_SPLIT 166 q330 q331
XSPLIT167 LSmitll_SPLIT 167 q332 q333
XSPLIT168 LSmitll_SPLIT 168 q334 q335
XSPLIT169 LSmitll_SPLIT 169 q336 q337
XSPLIT170 LSmitll_SPLIT 170 q338 q339
XSPLIT171 LSmitll_SPLIT 171 q340 q341
XSPLIT172 LSmitll_SPLIT 172 q342 q343
XSPLIT173 LSmitll_SPLIT 173 q344 q345
XSPLIT174 LSmitll_SPLIT 174 q346 q347
XSPLIT175 LSmitll_SPLIT 175 q348 q349
XSPLIT176 LSmitll_SPLIT 176 q350 q351
XSPLIT177 LSmitll_SPLIT 177 q352 q353
XSPLIT178 LSmitll_SPLIT 178 q354 q355
XSPLIT179 LSmitll_SPLIT 179 q356 q357
XSPLIT180 LSmitll_SPLIT 180 q358 q359
XSPLIT181 LSmitll_SPLIT 181 q360 q361
XSPLIT182 LSmitll_SPLIT 182 q362 q363
XSPLIT183 LSmitll_SPLIT 183 q364 q365
XSPLIT184 LSmitll_SPLIT 184 q366 q367
XSPLIT185 LSmitll_SPLIT 185 q368 q369
XSPLIT186 LSmitll_SPLIT 186 q370 q371
XSPLIT187 LSmitll_SPLIT 187 q372 q373
XSPLIT188 LSmitll_SPLIT 188 q374 q375
XSPLIT189 LSmitll_SPLIT 189 q376 q377
XSPLIT190 LSmitll_SPLIT 190 q378 q379
XSPLIT191 LSmitll_SPLIT 191 q380 q381
XSPLIT192 LSmitll_SPLIT 192 q382 q383
XSPLIT193 LSmitll_SPLIT 193 q384 q385
XSPLIT194 LSmitll_SPLIT 194 q386 q387
XSPLIT195 LSmitll_SPLIT 195 q388 q389
XSPLIT196 LSmitll_SPLIT 196 q390 q391
XSPLIT197 LSmitll_SPLIT 197 q392 q393
XSPLIT198 LSmitll_SPLIT 198 q394 q395
XSPLIT199 LSmitll_SPLIT 199 q396 q397
XSPLIT200 LSmitll_SPLIT 200 q398 q399
XSPLIT201 LSmitll_SPLIT 201 q400 q401
XSPLIT202 LSmitll_SPLIT 202 q402 q403
XSPLIT203 LSmitll_SPLIT 203 q404 q405
XSPLIT204 LSmitll_SPLIT 204 q406 q407
XSPLIT205 LSmitll_SPLIT 205 q408 q409
XSPLIT206 LSmitll_SPLIT 206 q410 q411
XSPLIT207 LSmitll_SPLIT 207 q412 q413
XSPLIT208 LSmitll_SPLIT 208 q414 q415
XSPLIT209 LSmitll_SPLIT 209 q416 q417
XSPLIT210 LSmitll_SPLIT 210 q418 q419
XSPLIT211 LSmitll_SPLIT 211 q420 q421
XSPLIT212 LSmitll_SPLIT 212 q422 q423
XSPLIT213 LSmitll_SPLIT 213 q424 q425
XSPLIT214 LSmitll_SPLIT 214 q426 q427
XSPLIT215 LSmitll_SPLIT 215 q428 q429
XSPLIT216 LSmitll_SPLIT 216 q430 q431
XSPLIT217 LSmitll_SPLIT 217 q432 q433
XSPLIT218 LSmitll_SPLIT 218 q434 q435
XSPLIT219 LSmitll_SPLIT 219 q436 q437
XSPLIT220 LSmitll_SPLIT 220 q438 q439
XSPLIT221 LSmitll_SPLIT 221 q440 q441
XSPLIT222 LSmitll_SPLIT 222 q442 q443
XSPLIT223 LSmitll_SPLIT 223 q444 q445
XSPLIT224 LSmitll_SPLIT 224 q446 q447
XSPLIT225 LSmitll_SPLIT 225 q448 q449
XSPLIT226 LSmitll_SPLIT 226 q450 q451
XSPLIT227 LSmitll_SPLIT 227 q452 q453
XSPLIT228 LSmitll_SPLIT 228 q454 q455
XSPLIT229 LSmitll_SPLIT 229 q456 q457
XSPLIT230 LSmitll_SPLIT 230 q458 q459
XSPLIT231 LSmitll_SPLIT 231 q460 q461
XSPLIT232 LSmitll_SPLIT 232 q462 q463
XSPLIT233 LSmitll_SPLIT 233 q464 q465
XSPLIT234 LSmitll_SPLIT 234 q466 q467
XSPLIT235 LSmitll_SPLIT 235 q468 q469
XSPLIT236 LSmitll_SPLIT 236 q470 q471
XSPLIT237 LSmitll_SPLIT 237 q472 q473
XSPLIT238 LSmitll_SPLIT 238 q474 q475
XSPLIT239 LSmitll_SPLIT 239 q476 q477
XSPLIT240 LSmitll_SPLIT 240 q478 q479
XSPLIT241 LSmitll_SPLIT 241 q480 q481
XSPLIT242 LSmitll_SPLIT 242 q482 q483
XSPLIT243 LSmitll_SPLIT 243 q484 q485
XSPLIT244 LSmitll_SPLIT 244 q486 q487
XSPLIT245 LSmitll_SPLIT 245 q488 q489
XSPLIT246 LSmitll_SPLIT 246 q490 q491
XSPLIT247 LSmitll_SPLIT 247 q492 q493
XSPLIT248 LSmitll_SPLIT 248 q494 q495
XSPLIT249 LSmitll_SPLIT 249 q496 q497
XSPLIT250 LSmitll_SPLIT 250 q498 q499
XSPLIT251 LSmitll_SPLIT 251 q500 q501
XSPLIT252 LSmitll_SPLIT 252 q502 q503
XSPLIT253 LSmitll_SPLIT 253 q504 q505
XSPLIT254 LSmitll_SPLIT 254 q506 q507
XSPLIT255 LSmitll_SPLIT 255 q508 q509
XSPLIT256 LSmitll_SPLIT 256 q510 q511
XSPLIT257 LSmitll_SPLIT 257 q512 q513
XSPLIT258 LSmitll_SPLIT 258 q514 q515
XSPLIT259 LSmitll_SPLIT 259 q516 q517
XSPLIT260 LSmitll_SPLIT 260 q518 q519
XSPLIT261 LSmitll_SPLIT 261 q520 q521
XSPLIT262 LSmitll_SPLIT 262 q522 q523
XSPLIT263 LSmitll_SPLIT 263 q524 q525
XSPLIT264 LSmitll_SPLIT 264 q526 q527
XSPLIT265 LSmitll_SPLIT 265 q528 q529
XSPLIT266 LSmitll_SPLIT 266 q530 q531
XSPLIT267 LSmitll_SPLIT 267 q532 q533
XSPLIT268 LSmitll_SPLIT 268 q534 q535
XSPLIT269 LSmitll_SPLIT 269 q536 q537
XSPLIT270 LSmitll_SPLIT 270 q538 q539
XSPLIT271 LSmitll_SPLIT 271 q540 q541
XSPLIT272 LSmitll_SPLIT 272 q542 q543
XSPLIT273 LSmitll_SPLIT 273 q544 q545
XSPLIT274 LSmitll_SPLIT 274 q546 q547
XSPLIT275 LSmitll_SPLIT 275 q548 q549
XSPLIT276 LSmitll_SPLIT 276 q550 q551
XSPLIT277 LSmitll_SPLIT 277 q552 q553
XSPLIT278 LSmitll_SPLIT 278 q554 q555
XSPLIT279 LSmitll_SPLIT 279 q556 q557
XSPLIT280 LSmitll_SPLIT 280 q558 q559
XSPLIT281 LSmitll_SPLIT 281 q560 q561
XSPLIT282 LSmitll_SPLIT 282 q562 q563
XSPLIT283 LSmitll_SPLIT 283 q564 q565
XSPLIT284 LSmitll_SPLIT 284 q566 q567
XSPLIT285 LSmitll_SPLIT 285 q568 q569
XSPLIT286 LSmitll_SPLIT 286 q570 q571
XSPLIT287 LSmitll_SPLIT 287 q572 q573
XSPLIT288 LSmitll_SPLIT 288 q574 q575
XSPLIT289 LSmitll_SPLIT 289 q576 q577
XSPLIT290 LSmitll_SPLIT 290 q578 q579
XSPLIT291 LSmitll_SPLIT 291 q580 q581
XSPLIT292 LSmitll_SPLIT 292 q582 q583
XSPLIT293 LSmitll_SPLIT 293 q584 q585
XSPLIT294 LSmitll_SPLIT 294 q586 q587
XSPLIT295 LSmitll_SPLIT 295 q588 q589
XSPLIT296 LSmitll_SPLIT 296 q590 q591
XSPLIT297 LSmitll_SPLIT 297 q592 q593
XSPLIT298 LSmitll_SPLIT 298 q594 q595
XSPLIT299 LSmitll_SPLIT 299 q596 q597
XSPLIT300 LSmitll_SPLIT 300 q598 q599
XSPLIT301 LSmitll_SPLIT 301 q600 q601
XSPLIT302 LSmitll_SPLIT 302 q602 q603
XSPLIT303 LSmitll_SPLIT 303 q604 q605
XSPLIT304 LSmitll_SPLIT 304 q606 q607
XSPLIT305 LSmitll_SPLIT 305 q608 q609
XSPLIT306 LSmitll_SPLIT 306 q610 q611
XSPLIT307 LSmitll_SPLIT 307 q612 q613
XSPLIT308 LSmitll_SPLIT 308 q614 q615
XSPLIT309 LSmitll_SPLIT 309 q616 q617
XSPLIT310 LSmitll_SPLIT 310 q618 q619
XSPLIT311 LSmitll_SPLIT 311 q620 q621
XSPLIT312 LSmitll_SPLIT 312 q622 q623
XSPLIT313 LSmitll_SPLIT 313 q624 q625
XSPLIT314 LSmitll_SPLIT 314 q626 q627
XSPLIT315 LSmitll_SPLIT 315 q628 q629
XSPLIT316 LSmitll_SPLIT 316 q630 q631
XSPLIT317 LSmitll_SPLIT 317 q632 q633
XSPLIT318 LSmitll_SPLIT 318 q634 q635
XSPLIT319 LSmitll_SPLIT 319 q636 q637
XSPLIT320 LSmitll_SPLIT 320 q638 q639
XSPLIT321 LSmitll_SPLIT 321 q640 q641
XSPLIT322 LSmitll_SPLIT 322 q642 q643
XSPLIT323 LSmitll_SPLIT 323 q644 q645
XSPLIT324 LSmitll_SPLIT 324 q646 q647
XSPLIT325 LSmitll_SPLIT 325 q648 q649
XSPLIT326 LSmitll_SPLIT 326 q650 q651
XSPLIT327 LSmitll_SPLIT 327 q652 q653
XSPLIT328 LSmitll_SPLIT 328 q654 q655
XSPLIT329 LSmitll_SPLIT 329 q656 q657
XSPLIT330 LSmitll_SPLIT 330 q658 q659
XSPLIT331 LSmitll_SPLIT 331 q660 q661
XSPLIT332 LSmitll_SPLIT 332 q662 q663
XSPLIT333 LSmitll_SPLIT 333 q664 q665
XSPLIT334 LSmitll_SPLIT 334 q666 q667
XSPLIT335 LSmitll_SPLIT 335 q668 q669
XSPLIT336 LSmitll_SPLIT 336 q670 q671
XSPLIT337 LSmitll_SPLIT 337 q672 q673
XSPLIT338 LSmitll_SPLIT 338 q674 q675
XSPLIT339 LSmitll_SPLIT 339 q676 q677
XSPLIT340 LSmitll_SPLIT 340 q678 q679
XSPLIT341 LSmitll_SPLIT 341 q680 q681
XSPLIT342 LSmitll_SPLIT 342 q682 q683
XSPLIT343 LSmitll_SPLIT 343 q684 q685
XSPLIT344 LSmitll_SPLIT 344 q686 q687
XSPLIT345 LSmitll_SPLIT 345 q688 q689
XSPLIT346 LSmitll_SPLIT 346 q690 q691
XSPLIT347 LSmitll_SPLIT 347 q692 q693
XSPLIT348 LSmitll_SPLIT 348 q694 q695
XSPLIT349 LSmitll_SPLIT 349 q696 q697
XSPLIT350 LSmitll_SPLIT 350 q698 q699
XSPLIT351 LSmitll_SPLIT 351 q700 q701
XSPLIT352 LSmitll_SPLIT 352 q702 q703
XSPLIT353 LSmitll_SPLIT 353 q704 q705
XSPLIT354 LSmitll_SPLIT 354 q706 q707
XSPLIT355 LSmitll_SPLIT 355 q708 q709
XSPLIT356 LSmitll_SPLIT 356 q710 q711
XSPLIT357 LSmitll_SPLIT 357 q712 q713
XSPLIT358 LSmitll_SPLIT 358 q714 q715
XSPLIT359 LSmitll_SPLIT 359 q716 q717
XSPLIT360 LSmitll_SPLIT 360 q718 q719
XSPLIT361 LSmitll_SPLIT 361 q720 q721
XSPLIT362 LSmitll_SPLIT 362 q722 q723
XSPLIT363 LSmitll_SPLIT 363 q724 q725
XSPLIT364 LSmitll_SPLIT 364 q726 q727
XSPLIT365 LSmitll_SPLIT 365 q728 q729
XSPLIT366 LSmitll_SPLIT 366 q730 q731
XSPLIT367 LSmitll_SPLIT 367 q732 q733
XSPLIT368 LSmitll_SPLIT 368 q734 q735
XSPLIT369 LSmitll_SPLIT 369 q736 q737
XSPLIT370 LSmitll_SPLIT 370 q738 q739
XSPLIT371 LSmitll_SPLIT 371 q740 q741
XSPLIT372 LSmitll_SPLIT 372 q742 q743
XSPLIT373 LSmitll_SPLIT 373 q744 q745
XSPLIT374 LSmitll_SPLIT 374 q746 q747
XSPLIT375 LSmitll_SPLIT 375 q748 q749
XSPLIT376 LSmitll_SPLIT 376 q750 q751
XSPLIT377 LSmitll_SPLIT 377 q752 q753
XSPLIT378 LSmitll_SPLIT 378 q754 q755
XSPLIT379 LSmitll_SPLIT 379 q756 q757
XSPLIT380 LSmitll_SPLIT 380 q758 q759
XSPLIT381 LSmitll_SPLIT 381 q760 q761
XSPLIT382 LSmitll_SPLIT 382 q762 q763
XSPLIT383 LSmitll_SPLIT 383 q764 q765
XSPLIT384 LSmitll_SPLIT 384 q766 q767
XSPLIT385 LSmitll_SPLIT 385 q768 q769
XSPLIT386 LSmitll_SPLIT 386 q770 q771
XSPLIT387 LSmitll_SPLIT 387 q772 q773
XSPLIT388 LSmitll_SPLIT 388 q774 q775
XSPLIT389 LSmitll_SPLIT 389 q776 q777
XSPLIT390 LSmitll_SPLIT 390 q778 q779
XSPLIT391 LSmitll_SPLIT 391 q780 q781
XSPLIT392 LSmitll_SPLIT 392 q782 q783
XSPLIT393 LSmitll_SPLIT 393 q784 q785
XSPLIT394 LSmitll_SPLIT 394 q786 q787
XSPLIT395 LSmitll_SPLIT 395 q788 q789
XSPLIT396 LSmitll_SPLIT 396 q790 q791
XSPLIT397 LSmitll_SPLIT 397 q792 q793
XSPLIT398 LSmitll_SPLIT 398 q794 q795
XSPLIT399 LSmitll_SPLIT 399 q796 q797
XSPLIT400 LSmitll_SPLIT 400 q798 q799
XSPLIT401 LSmitll_SPLIT 401 q800 q801
XSPLIT402 LSmitll_SPLIT 402 q802 q803
XSPLIT403 LSmitll_SPLIT 403 q804 q805
XSPLIT404 LSmitll_SPLIT 404 q806 q807
XSPLIT405 LSmitll_SPLIT 405 q808 q809
XSPLIT406 LSmitll_SPLIT 406 q810 q811
XSPLIT407 LSmitll_SPLIT 407 q812 q813
XSPLIT408 LSmitll_SPLIT 408 q814 q815
XSPLIT409 LSmitll_SPLIT 409 q816 q817
XSPLIT410 LSmitll_SPLIT 410 q818 q819
XSPLIT411 LSmitll_SPLIT 411 q820 q821
XSPLIT412 LSmitll_SPLIT 412 q822 q823
XSPLIT413 LSmitll_SPLIT 413 q824 q825
XSPLIT414 LSmitll_SPLIT 414 q826 q827
XSPLIT415 LSmitll_SPLIT 415 q828 q829
XSPLIT416 LSmitll_SPLIT 416 q830 q831
XSPLIT417 LSmitll_SPLIT 417 q832 q833
XSPLIT418 LSmitll_SPLIT 418 q834 q835
XSPLIT419 LSmitll_SPLIT 419 q836 q837
XSPLIT420 LSmitll_SPLIT 420 q838 q839
XSPLIT421 LSmitll_SPLIT 421 q840 q841
XSPLIT422 LSmitll_SPLIT 422 q842 q843
XSPLIT423 LSmitll_SPLIT 423 q844 q845
XSPLIT424 LSmitll_SPLIT 424 q846 q847
.ends 1_to_848_split
* change up

.subckt 1_to_1024_split a q0 q1 q2 q3 q4 q5 q6 q7 q8 q9 q10 q11 q12 q13 q14 q15 q16 q17 q18 q19 q20 q21 q22 q23 q24 q25 q26 q27 q28 q29 q30 q31 q32 q33 q34 q35 q36 q37 q38 q39 q40 q41 q42 q43 q44 q45 q46 q47 q48 q49 q50 q51 q52 q53 q54 q55 q56 q57 q58 q59 q60 q61 q62 q63 q64 q65 q66 q67 q68 q69 q70 q71 q72 q73 q74 q75 q76 q77 q78 q79 q80 q81 q82 q83 q84 q85 q86 q87 q88 q89 q90 q91 q92 q93 q94 q95 q96 q97 q98 q99 q100 q101 q102 q103 q104 q105 q106 q107 q108 q109 q110 q111 q112 q113 q114 q115 q116 q117 q118 q119 q120 q121 q122 q123 q124 q125 q126 q127 q128 q129 q130 q131 q132 q133 q134 q135 q136 q137 q138 q139 q140 q141 q142 q143 q144 q145 q146 q147 q148 q149 q150 q151 q152 q153 q154 q155 q156 q157 q158 q159 q160 q161 q162 q163 q164 q165 q166 q167 q168 q169 q170 q171 q172 q173 q174 q175 q176 q177 q178 q179 q180 q181 q182 q183 q184 q185 q186 q187 q188 q189 q190 q191 q192 q193 q194 q195 q196 q197 q198 q199 q200 q201 q202 q203 q204 q205 q206 q207 q208 q209 q210 q211 q212 q213 q214 q215 q216 q217 q218 q219 q220 q221 q222 q223 q224 q225 q226 q227 q228 q229 q230 q231 q232 q233 q234 q235 q236 q237 q238 q239 q240 q241 q242 q243 q244 q245 q246 q247 q248 q249 q250 q251 q252 q253 q254 q255 q256 q257 q258 q259 q260 q261 q262 q263 q264 q265 q266 q267 q268 q269 q270 q271 q272 q273 q274 q275 q276 q277 q278 q279 q280 q281 q282 q283 q284 q285 q286 q287 q288 q289 q290 q291 q292 q293 q294 q295 q296 q297 q298 q299 q300 q301 q302 q303 q304 q305 q306 q307 q308 q309 q310 q311 q312 q313 q314 q315 q316 q317 q318 q319 q320 q321 q322 q323 q324 q325 q326 q327 q328 q329 q330 q331 q332 q333 q334 q335 q336 q337 q338 q339 q340 q341 q342 q343 q344 q345 q346 q347 q348 q349 q350 q351 q352 q353 q354 q355 q356 q357 q358 q359 q360 q361 q362 q363 q364 q365 q366 q367 q368 q369 q370 q371 q372 q373 q374 q375 q376 q377 q378 q379 q380 q381 q382 q383 q384 q385 q386 q387 q388 q389 q390 q391 q392 q393 q394 q395 q396 q397 q398 q399 q400 q401 q402 q403 q404 q405 q406 q407 q408 q409 q410 q411 q412 q413 q414 q415 q416 q417 q418 q419 q420 q421 q422 q423 q424 q425 q426 q427 q428 q429 q430 q431 q432 q433 q434 q435 q436 q437 q438 q439 q440 q441 q442 q443 q444 q445 q446 q447 q448 q449 q450 q451 q452 q453 q454 q455 q456 q457 q458 q459 q460 q461 q462 q463 q464 q465 q466 q467 q468 q469 q470 q471 q472 q473 q474 q475 q476 q477 q478 q479 q480 q481 q482 q483 q484 q485 q486 q487 q488 q489 q490 q491 q492 q493 q494 q495 q496 q497 q498 q499 q500 q501 q502 q503 q504 q505 q506 q507 q508 q509 q510 q511 q512 q513 q514 q515 q516 q517 q518 q519 q520 q521 q522 q523 q524 q525 q526 q527 q528 q529 q530 q531 q532 q533 q534 q535 q536 q537 q538 q539 q540 q541 q542 q543 q544 q545 q546 q547 q548 q549 q550 q551 q552 q553 q554 q555 q556 q557 q558 q559 q560 q561 q562 q563 q564 q565 q566 q567 q568 q569 q570 q571 q572 q573 q574 q575 q576 q577 q578 q579 q580 q581 q582 q583 q584 q585 q586 q587 q588 q589 q590 q591 q592 q593 q594 q595 q596 q597 q598 q599 q600 q601 q602 q603 q604 q605 q606 q607 q608 q609 q610 q611 q612 q613 q614 q615 q616 q617 q618 q619 q620 q621 q622 q623 q624 q625 q626 q627 q628 q629 q630 q631 q632 q633 q634 q635 q636 q637 q638 q639 q640 q641 q642 q643 q644 q645 q646 q647 q648 q649 q650 q651 q652 q653 q654 q655 q656 q657 q658 q659 q660 q661 q662 q663 q664 q665 q666 q667 q668 q669 q670 q671 q672 q673 q674 q675 q676 q677 q678 q679 q680 q681 q682 q683 q684 q685 q686 q687 q688 q689 q690 q691 q692 q693 q694 q695 q696 q697 q698 q699 q700 q701 q702 q703 q704 q705 q706 q707 q708 q709 q710 q711 q712 q713 q714 q715 q716 q717 q718 q719 q720 q721 q722 q723 q724 q725 q726 q727 q728 q729 q730 q731 q732 q733 q734 q735 q736 q737 q738 q739 q740 q741 q742 q743 q744 q745 q746 q747 q748 q749 q750 q751 q752 q753 q754 q755 q756 q757 q758 q759 q760 q761 q762 q763 q764 q765 q766 q767 q768 q769 q770 q771 q772 q773 q774 q775 q776 q777 q778 q779 q780 q781 q782 q783 q784 q785 q786 q787 q788 q789 q790 q791 q792 q793 q794 q795 q796 q797 q798 q799 q800 q801 q802 q803 q804 q805 q806 q807 q808 q809 q810 q811 q812 q813 q814 q815 q816 q817 q818 q819 q820 q821 q822 q823 q824 q825 q826 q827 q828 q829 q830 q831 q832 q833 q834 q835 q836 q837 q838 q839 q840 q841 q842 q843 q844 q845 q846 q847 q848 q849 q850 q851 q852 q853 q854 q855 q856 q857 q858 q859 q860 q861 q862 q863 q864 q865 q866 q867 q868 q869 q870 q871 q872 q873 q874 q875 q876 q877 q878 q879 q880 q881 q882 q883 q884 q885 q886 q887 q888 q889 q890 q891 q892 q893 q894 q895 q896 q897 q898 q899 q900 q901 q902 q903 q904 q905 q906 q907 q908 q909 q910 q911 q912 q913 q914 q915 q916 q917 q918 q919 q920 q921 q922 q923 q924 q925 q926 q927 q928 q929 q930 q931 q932 q933 q934 q935 q936 q937 q938 q939 q940 q941 q942 q943 q944 q945 q946 q947 q948 q949 q950 q951 q952 q953 q954 q955 q956 q957 q958 q959 q960 q961 q962 q963 q964 q965 q966 q967 q968 q969 q970 q971 q972 q973 q974 q975 q976 q977 q978 q979 q980 q981 q982 q983 q984 q985 q986 q987 q988 q989 q990 q991 q992 q993 q994 q995 q996 q997 q998 q999 q1000 q1001 q1002 q1003 q1004 q1005 q1006 q1007 q1008 q1009 q1010 q1011 q1012 q1013 q1014 q1015 q1016 q1017 q1018 q1019 q1020 q1021 q1022 q1023 
XSPLIT_512 1_to_512_split a 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510 511 512 
XSPLIT1 LSmitll_SPLIT 1 q0 q1
XSPLIT2 LSmitll_SPLIT 2 q2 q3
XSPLIT3 LSmitll_SPLIT 3 q4 q5
XSPLIT4 LSmitll_SPLIT 4 q6 q7
XSPLIT5 LSmitll_SPLIT 5 q8 q9
XSPLIT6 LSmitll_SPLIT 6 q10 q11
XSPLIT7 LSmitll_SPLIT 7 q12 q13
XSPLIT8 LSmitll_SPLIT 8 q14 q15
XSPLIT9 LSmitll_SPLIT 9 q16 q17
XSPLIT10 LSmitll_SPLIT 10 q18 q19
XSPLIT11 LSmitll_SPLIT 11 q20 q21
XSPLIT12 LSmitll_SPLIT 12 q22 q23
XSPLIT13 LSmitll_SPLIT 13 q24 q25
XSPLIT14 LSmitll_SPLIT 14 q26 q27
XSPLIT15 LSmitll_SPLIT 15 q28 q29
XSPLIT16 LSmitll_SPLIT 16 q30 q31
XSPLIT17 LSmitll_SPLIT 17 q32 q33
XSPLIT18 LSmitll_SPLIT 18 q34 q35
XSPLIT19 LSmitll_SPLIT 19 q36 q37
XSPLIT20 LSmitll_SPLIT 20 q38 q39
XSPLIT21 LSmitll_SPLIT 21 q40 q41
XSPLIT22 LSmitll_SPLIT 22 q42 q43
XSPLIT23 LSmitll_SPLIT 23 q44 q45
XSPLIT24 LSmitll_SPLIT 24 q46 q47
XSPLIT25 LSmitll_SPLIT 25 q48 q49
XSPLIT26 LSmitll_SPLIT 26 q50 q51
XSPLIT27 LSmitll_SPLIT 27 q52 q53
XSPLIT28 LSmitll_SPLIT 28 q54 q55
XSPLIT29 LSmitll_SPLIT 29 q56 q57
XSPLIT30 LSmitll_SPLIT 30 q58 q59
XSPLIT31 LSmitll_SPLIT 31 q60 q61
XSPLIT32 LSmitll_SPLIT 32 q62 q63
XSPLIT33 LSmitll_SPLIT 33 q64 q65
XSPLIT34 LSmitll_SPLIT 34 q66 q67
XSPLIT35 LSmitll_SPLIT 35 q68 q69
XSPLIT36 LSmitll_SPLIT 36 q70 q71
XSPLIT37 LSmitll_SPLIT 37 q72 q73
XSPLIT38 LSmitll_SPLIT 38 q74 q75
XSPLIT39 LSmitll_SPLIT 39 q76 q77
XSPLIT40 LSmitll_SPLIT 40 q78 q79
XSPLIT41 LSmitll_SPLIT 41 q80 q81
XSPLIT42 LSmitll_SPLIT 42 q82 q83
XSPLIT43 LSmitll_SPLIT 43 q84 q85
XSPLIT44 LSmitll_SPLIT 44 q86 q87
XSPLIT45 LSmitll_SPLIT 45 q88 q89
XSPLIT46 LSmitll_SPLIT 46 q90 q91
XSPLIT47 LSmitll_SPLIT 47 q92 q93
XSPLIT48 LSmitll_SPLIT 48 q94 q95
XSPLIT49 LSmitll_SPLIT 49 q96 q97
XSPLIT50 LSmitll_SPLIT 50 q98 q99
XSPLIT51 LSmitll_SPLIT 51 q100 q101
XSPLIT52 LSmitll_SPLIT 52 q102 q103
XSPLIT53 LSmitll_SPLIT 53 q104 q105
XSPLIT54 LSmitll_SPLIT 54 q106 q107
XSPLIT55 LSmitll_SPLIT 55 q108 q109
XSPLIT56 LSmitll_SPLIT 56 q110 q111
XSPLIT57 LSmitll_SPLIT 57 q112 q113
XSPLIT58 LSmitll_SPLIT 58 q114 q115
XSPLIT59 LSmitll_SPLIT 59 q116 q117
XSPLIT60 LSmitll_SPLIT 60 q118 q119
XSPLIT61 LSmitll_SPLIT 61 q120 q121
XSPLIT62 LSmitll_SPLIT 62 q122 q123
XSPLIT63 LSmitll_SPLIT 63 q124 q125
XSPLIT64 LSmitll_SPLIT 64 q126 q127
XSPLIT65 LSmitll_SPLIT 65 q128 q129
XSPLIT66 LSmitll_SPLIT 66 q130 q131
XSPLIT67 LSmitll_SPLIT 67 q132 q133
XSPLIT68 LSmitll_SPLIT 68 q134 q135
XSPLIT69 LSmitll_SPLIT 69 q136 q137
XSPLIT70 LSmitll_SPLIT 70 q138 q139
XSPLIT71 LSmitll_SPLIT 71 q140 q141
XSPLIT72 LSmitll_SPLIT 72 q142 q143
XSPLIT73 LSmitll_SPLIT 73 q144 q145
XSPLIT74 LSmitll_SPLIT 74 q146 q147
XSPLIT75 LSmitll_SPLIT 75 q148 q149
XSPLIT76 LSmitll_SPLIT 76 q150 q151
XSPLIT77 LSmitll_SPLIT 77 q152 q153
XSPLIT78 LSmitll_SPLIT 78 q154 q155
XSPLIT79 LSmitll_SPLIT 79 q156 q157
XSPLIT80 LSmitll_SPLIT 80 q158 q159
XSPLIT81 LSmitll_SPLIT 81 q160 q161
XSPLIT82 LSmitll_SPLIT 82 q162 q163
XSPLIT83 LSmitll_SPLIT 83 q164 q165
XSPLIT84 LSmitll_SPLIT 84 q166 q167
XSPLIT85 LSmitll_SPLIT 85 q168 q169
XSPLIT86 LSmitll_SPLIT 86 q170 q171
XSPLIT87 LSmitll_SPLIT 87 q172 q173
XSPLIT88 LSmitll_SPLIT 88 q174 q175
XSPLIT89 LSmitll_SPLIT 89 q176 q177
XSPLIT90 LSmitll_SPLIT 90 q178 q179
XSPLIT91 LSmitll_SPLIT 91 q180 q181
XSPLIT92 LSmitll_SPLIT 92 q182 q183
XSPLIT93 LSmitll_SPLIT 93 q184 q185
XSPLIT94 LSmitll_SPLIT 94 q186 q187
XSPLIT95 LSmitll_SPLIT 95 q188 q189
XSPLIT96 LSmitll_SPLIT 96 q190 q191
XSPLIT97 LSmitll_SPLIT 97 q192 q193
XSPLIT98 LSmitll_SPLIT 98 q194 q195
XSPLIT99 LSmitll_SPLIT 99 q196 q197
XSPLIT100 LSmitll_SPLIT 100 q198 q199
XSPLIT101 LSmitll_SPLIT 101 q200 q201
XSPLIT102 LSmitll_SPLIT 102 q202 q203
XSPLIT103 LSmitll_SPLIT 103 q204 q205
XSPLIT104 LSmitll_SPLIT 104 q206 q207
XSPLIT105 LSmitll_SPLIT 105 q208 q209
XSPLIT106 LSmitll_SPLIT 106 q210 q211
XSPLIT107 LSmitll_SPLIT 107 q212 q213
XSPLIT108 LSmitll_SPLIT 108 q214 q215
XSPLIT109 LSmitll_SPLIT 109 q216 q217
XSPLIT110 LSmitll_SPLIT 110 q218 q219
XSPLIT111 LSmitll_SPLIT 111 q220 q221
XSPLIT112 LSmitll_SPLIT 112 q222 q223
XSPLIT113 LSmitll_SPLIT 113 q224 q225
XSPLIT114 LSmitll_SPLIT 114 q226 q227
XSPLIT115 LSmitll_SPLIT 115 q228 q229
XSPLIT116 LSmitll_SPLIT 116 q230 q231
XSPLIT117 LSmitll_SPLIT 117 q232 q233
XSPLIT118 LSmitll_SPLIT 118 q234 q235
XSPLIT119 LSmitll_SPLIT 119 q236 q237
XSPLIT120 LSmitll_SPLIT 120 q238 q239
XSPLIT121 LSmitll_SPLIT 121 q240 q241
XSPLIT122 LSmitll_SPLIT 122 q242 q243
XSPLIT123 LSmitll_SPLIT 123 q244 q245
XSPLIT124 LSmitll_SPLIT 124 q246 q247
XSPLIT125 LSmitll_SPLIT 125 q248 q249
XSPLIT126 LSmitll_SPLIT 126 q250 q251
XSPLIT127 LSmitll_SPLIT 127 q252 q253
XSPLIT128 LSmitll_SPLIT 128 q254 q255
XSPLIT129 LSmitll_SPLIT 129 q256 q257
XSPLIT130 LSmitll_SPLIT 130 q258 q259
XSPLIT131 LSmitll_SPLIT 131 q260 q261
XSPLIT132 LSmitll_SPLIT 132 q262 q263
XSPLIT133 LSmitll_SPLIT 133 q264 q265
XSPLIT134 LSmitll_SPLIT 134 q266 q267
XSPLIT135 LSmitll_SPLIT 135 q268 q269
XSPLIT136 LSmitll_SPLIT 136 q270 q271
XSPLIT137 LSmitll_SPLIT 137 q272 q273
XSPLIT138 LSmitll_SPLIT 138 q274 q275
XSPLIT139 LSmitll_SPLIT 139 q276 q277
XSPLIT140 LSmitll_SPLIT 140 q278 q279
XSPLIT141 LSmitll_SPLIT 141 q280 q281
XSPLIT142 LSmitll_SPLIT 142 q282 q283
XSPLIT143 LSmitll_SPLIT 143 q284 q285
XSPLIT144 LSmitll_SPLIT 144 q286 q287
XSPLIT145 LSmitll_SPLIT 145 q288 q289
XSPLIT146 LSmitll_SPLIT 146 q290 q291
XSPLIT147 LSmitll_SPLIT 147 q292 q293
XSPLIT148 LSmitll_SPLIT 148 q294 q295
XSPLIT149 LSmitll_SPLIT 149 q296 q297
XSPLIT150 LSmitll_SPLIT 150 q298 q299
XSPLIT151 LSmitll_SPLIT 151 q300 q301
XSPLIT152 LSmitll_SPLIT 152 q302 q303
XSPLIT153 LSmitll_SPLIT 153 q304 q305
XSPLIT154 LSmitll_SPLIT 154 q306 q307
XSPLIT155 LSmitll_SPLIT 155 q308 q309
XSPLIT156 LSmitll_SPLIT 156 q310 q311
XSPLIT157 LSmitll_SPLIT 157 q312 q313
XSPLIT158 LSmitll_SPLIT 158 q314 q315
XSPLIT159 LSmitll_SPLIT 159 q316 q317
XSPLIT160 LSmitll_SPLIT 160 q318 q319
XSPLIT161 LSmitll_SPLIT 161 q320 q321
XSPLIT162 LSmitll_SPLIT 162 q322 q323
XSPLIT163 LSmitll_SPLIT 163 q324 q325
XSPLIT164 LSmitll_SPLIT 164 q326 q327
XSPLIT165 LSmitll_SPLIT 165 q328 q329
XSPLIT166 LSmitll_SPLIT 166 q330 q331
XSPLIT167 LSmitll_SPLIT 167 q332 q333
XSPLIT168 LSmitll_SPLIT 168 q334 q335
XSPLIT169 LSmitll_SPLIT 169 q336 q337
XSPLIT170 LSmitll_SPLIT 170 q338 q339
XSPLIT171 LSmitll_SPLIT 171 q340 q341
XSPLIT172 LSmitll_SPLIT 172 q342 q343
XSPLIT173 LSmitll_SPLIT 173 q344 q345
XSPLIT174 LSmitll_SPLIT 174 q346 q347
XSPLIT175 LSmitll_SPLIT 175 q348 q349
XSPLIT176 LSmitll_SPLIT 176 q350 q351
XSPLIT177 LSmitll_SPLIT 177 q352 q353
XSPLIT178 LSmitll_SPLIT 178 q354 q355
XSPLIT179 LSmitll_SPLIT 179 q356 q357
XSPLIT180 LSmitll_SPLIT 180 q358 q359
XSPLIT181 LSmitll_SPLIT 181 q360 q361
XSPLIT182 LSmitll_SPLIT 182 q362 q363
XSPLIT183 LSmitll_SPLIT 183 q364 q365
XSPLIT184 LSmitll_SPLIT 184 q366 q367
XSPLIT185 LSmitll_SPLIT 185 q368 q369
XSPLIT186 LSmitll_SPLIT 186 q370 q371
XSPLIT187 LSmitll_SPLIT 187 q372 q373
XSPLIT188 LSmitll_SPLIT 188 q374 q375
XSPLIT189 LSmitll_SPLIT 189 q376 q377
XSPLIT190 LSmitll_SPLIT 190 q378 q379
XSPLIT191 LSmitll_SPLIT 191 q380 q381
XSPLIT192 LSmitll_SPLIT 192 q382 q383
XSPLIT193 LSmitll_SPLIT 193 q384 q385
XSPLIT194 LSmitll_SPLIT 194 q386 q387
XSPLIT195 LSmitll_SPLIT 195 q388 q389
XSPLIT196 LSmitll_SPLIT 196 q390 q391
XSPLIT197 LSmitll_SPLIT 197 q392 q393
XSPLIT198 LSmitll_SPLIT 198 q394 q395
XSPLIT199 LSmitll_SPLIT 199 q396 q397
XSPLIT200 LSmitll_SPLIT 200 q398 q399
XSPLIT201 LSmitll_SPLIT 201 q400 q401
XSPLIT202 LSmitll_SPLIT 202 q402 q403
XSPLIT203 LSmitll_SPLIT 203 q404 q405
XSPLIT204 LSmitll_SPLIT 204 q406 q407
XSPLIT205 LSmitll_SPLIT 205 q408 q409
XSPLIT206 LSmitll_SPLIT 206 q410 q411
XSPLIT207 LSmitll_SPLIT 207 q412 q413
XSPLIT208 LSmitll_SPLIT 208 q414 q415
XSPLIT209 LSmitll_SPLIT 209 q416 q417
XSPLIT210 LSmitll_SPLIT 210 q418 q419
XSPLIT211 LSmitll_SPLIT 211 q420 q421
XSPLIT212 LSmitll_SPLIT 212 q422 q423
XSPLIT213 LSmitll_SPLIT 213 q424 q425
XSPLIT214 LSmitll_SPLIT 214 q426 q427
XSPLIT215 LSmitll_SPLIT 215 q428 q429
XSPLIT216 LSmitll_SPLIT 216 q430 q431
XSPLIT217 LSmitll_SPLIT 217 q432 q433
XSPLIT218 LSmitll_SPLIT 218 q434 q435
XSPLIT219 LSmitll_SPLIT 219 q436 q437
XSPLIT220 LSmitll_SPLIT 220 q438 q439
XSPLIT221 LSmitll_SPLIT 221 q440 q441
XSPLIT222 LSmitll_SPLIT 222 q442 q443
XSPLIT223 LSmitll_SPLIT 223 q444 q445
XSPLIT224 LSmitll_SPLIT 224 q446 q447
XSPLIT225 LSmitll_SPLIT 225 q448 q449
XSPLIT226 LSmitll_SPLIT 226 q450 q451
XSPLIT227 LSmitll_SPLIT 227 q452 q453
XSPLIT228 LSmitll_SPLIT 228 q454 q455
XSPLIT229 LSmitll_SPLIT 229 q456 q457
XSPLIT230 LSmitll_SPLIT 230 q458 q459
XSPLIT231 LSmitll_SPLIT 231 q460 q461
XSPLIT232 LSmitll_SPLIT 232 q462 q463
XSPLIT233 LSmitll_SPLIT 233 q464 q465
XSPLIT234 LSmitll_SPLIT 234 q466 q467
XSPLIT235 LSmitll_SPLIT 235 q468 q469
XSPLIT236 LSmitll_SPLIT 236 q470 q471
XSPLIT237 LSmitll_SPLIT 237 q472 q473
XSPLIT238 LSmitll_SPLIT 238 q474 q475
XSPLIT239 LSmitll_SPLIT 239 q476 q477
XSPLIT240 LSmitll_SPLIT 240 q478 q479
XSPLIT241 LSmitll_SPLIT 241 q480 q481
XSPLIT242 LSmitll_SPLIT 242 q482 q483
XSPLIT243 LSmitll_SPLIT 243 q484 q485
XSPLIT244 LSmitll_SPLIT 244 q486 q487
XSPLIT245 LSmitll_SPLIT 245 q488 q489
XSPLIT246 LSmitll_SPLIT 246 q490 q491
XSPLIT247 LSmitll_SPLIT 247 q492 q493
XSPLIT248 LSmitll_SPLIT 248 q494 q495
XSPLIT249 LSmitll_SPLIT 249 q496 q497
XSPLIT250 LSmitll_SPLIT 250 q498 q499
XSPLIT251 LSmitll_SPLIT 251 q500 q501
XSPLIT252 LSmitll_SPLIT 252 q502 q503
XSPLIT253 LSmitll_SPLIT 253 q504 q505
XSPLIT254 LSmitll_SPLIT 254 q506 q507
XSPLIT255 LSmitll_SPLIT 255 q508 q509
XSPLIT256 LSmitll_SPLIT 256 q510 q511
XSPLIT257 LSmitll_SPLIT 257 q512 q513
XSPLIT258 LSmitll_SPLIT 258 q514 q515
XSPLIT259 LSmitll_SPLIT 259 q516 q517
XSPLIT260 LSmitll_SPLIT 260 q518 q519
XSPLIT261 LSmitll_SPLIT 261 q520 q521
XSPLIT262 LSmitll_SPLIT 262 q522 q523
XSPLIT263 LSmitll_SPLIT 263 q524 q525
XSPLIT264 LSmitll_SPLIT 264 q526 q527
XSPLIT265 LSmitll_SPLIT 265 q528 q529
XSPLIT266 LSmitll_SPLIT 266 q530 q531
XSPLIT267 LSmitll_SPLIT 267 q532 q533
XSPLIT268 LSmitll_SPLIT 268 q534 q535
XSPLIT269 LSmitll_SPLIT 269 q536 q537
XSPLIT270 LSmitll_SPLIT 270 q538 q539
XSPLIT271 LSmitll_SPLIT 271 q540 q541
XSPLIT272 LSmitll_SPLIT 272 q542 q543
XSPLIT273 LSmitll_SPLIT 273 q544 q545
XSPLIT274 LSmitll_SPLIT 274 q546 q547
XSPLIT275 LSmitll_SPLIT 275 q548 q549
XSPLIT276 LSmitll_SPLIT 276 q550 q551
XSPLIT277 LSmitll_SPLIT 277 q552 q553
XSPLIT278 LSmitll_SPLIT 278 q554 q555
XSPLIT279 LSmitll_SPLIT 279 q556 q557
XSPLIT280 LSmitll_SPLIT 280 q558 q559
XSPLIT281 LSmitll_SPLIT 281 q560 q561
XSPLIT282 LSmitll_SPLIT 282 q562 q563
XSPLIT283 LSmitll_SPLIT 283 q564 q565
XSPLIT284 LSmitll_SPLIT 284 q566 q567
XSPLIT285 LSmitll_SPLIT 285 q568 q569
XSPLIT286 LSmitll_SPLIT 286 q570 q571
XSPLIT287 LSmitll_SPLIT 287 q572 q573
XSPLIT288 LSmitll_SPLIT 288 q574 q575
XSPLIT289 LSmitll_SPLIT 289 q576 q577
XSPLIT290 LSmitll_SPLIT 290 q578 q579
XSPLIT291 LSmitll_SPLIT 291 q580 q581
XSPLIT292 LSmitll_SPLIT 292 q582 q583
XSPLIT293 LSmitll_SPLIT 293 q584 q585
XSPLIT294 LSmitll_SPLIT 294 q586 q587
XSPLIT295 LSmitll_SPLIT 295 q588 q589
XSPLIT296 LSmitll_SPLIT 296 q590 q591
XSPLIT297 LSmitll_SPLIT 297 q592 q593
XSPLIT298 LSmitll_SPLIT 298 q594 q595
XSPLIT299 LSmitll_SPLIT 299 q596 q597
XSPLIT300 LSmitll_SPLIT 300 q598 q599
XSPLIT301 LSmitll_SPLIT 301 q600 q601
XSPLIT302 LSmitll_SPLIT 302 q602 q603
XSPLIT303 LSmitll_SPLIT 303 q604 q605
XSPLIT304 LSmitll_SPLIT 304 q606 q607
XSPLIT305 LSmitll_SPLIT 305 q608 q609
XSPLIT306 LSmitll_SPLIT 306 q610 q611
XSPLIT307 LSmitll_SPLIT 307 q612 q613
XSPLIT308 LSmitll_SPLIT 308 q614 q615
XSPLIT309 LSmitll_SPLIT 309 q616 q617
XSPLIT310 LSmitll_SPLIT 310 q618 q619
XSPLIT311 LSmitll_SPLIT 311 q620 q621
XSPLIT312 LSmitll_SPLIT 312 q622 q623
XSPLIT313 LSmitll_SPLIT 313 q624 q625
XSPLIT314 LSmitll_SPLIT 314 q626 q627
XSPLIT315 LSmitll_SPLIT 315 q628 q629
XSPLIT316 LSmitll_SPLIT 316 q630 q631
XSPLIT317 LSmitll_SPLIT 317 q632 q633
XSPLIT318 LSmitll_SPLIT 318 q634 q635
XSPLIT319 LSmitll_SPLIT 319 q636 q637
XSPLIT320 LSmitll_SPLIT 320 q638 q639
XSPLIT321 LSmitll_SPLIT 321 q640 q641
XSPLIT322 LSmitll_SPLIT 322 q642 q643
XSPLIT323 LSmitll_SPLIT 323 q644 q645
XSPLIT324 LSmitll_SPLIT 324 q646 q647
XSPLIT325 LSmitll_SPLIT 325 q648 q649
XSPLIT326 LSmitll_SPLIT 326 q650 q651
XSPLIT327 LSmitll_SPLIT 327 q652 q653
XSPLIT328 LSmitll_SPLIT 328 q654 q655
XSPLIT329 LSmitll_SPLIT 329 q656 q657
XSPLIT330 LSmitll_SPLIT 330 q658 q659
XSPLIT331 LSmitll_SPLIT 331 q660 q661
XSPLIT332 LSmitll_SPLIT 332 q662 q663
XSPLIT333 LSmitll_SPLIT 333 q664 q665
XSPLIT334 LSmitll_SPLIT 334 q666 q667
XSPLIT335 LSmitll_SPLIT 335 q668 q669
XSPLIT336 LSmitll_SPLIT 336 q670 q671
XSPLIT337 LSmitll_SPLIT 337 q672 q673
XSPLIT338 LSmitll_SPLIT 338 q674 q675
XSPLIT339 LSmitll_SPLIT 339 q676 q677
XSPLIT340 LSmitll_SPLIT 340 q678 q679
XSPLIT341 LSmitll_SPLIT 341 q680 q681
XSPLIT342 LSmitll_SPLIT 342 q682 q683
XSPLIT343 LSmitll_SPLIT 343 q684 q685
XSPLIT344 LSmitll_SPLIT 344 q686 q687
XSPLIT345 LSmitll_SPLIT 345 q688 q689
XSPLIT346 LSmitll_SPLIT 346 q690 q691
XSPLIT347 LSmitll_SPLIT 347 q692 q693
XSPLIT348 LSmitll_SPLIT 348 q694 q695
XSPLIT349 LSmitll_SPLIT 349 q696 q697
XSPLIT350 LSmitll_SPLIT 350 q698 q699
XSPLIT351 LSmitll_SPLIT 351 q700 q701
XSPLIT352 LSmitll_SPLIT 352 q702 q703
XSPLIT353 LSmitll_SPLIT 353 q704 q705
XSPLIT354 LSmitll_SPLIT 354 q706 q707
XSPLIT355 LSmitll_SPLIT 355 q708 q709
XSPLIT356 LSmitll_SPLIT 356 q710 q711
XSPLIT357 LSmitll_SPLIT 357 q712 q713
XSPLIT358 LSmitll_SPLIT 358 q714 q715
XSPLIT359 LSmitll_SPLIT 359 q716 q717
XSPLIT360 LSmitll_SPLIT 360 q718 q719
XSPLIT361 LSmitll_SPLIT 361 q720 q721
XSPLIT362 LSmitll_SPLIT 362 q722 q723
XSPLIT363 LSmitll_SPLIT 363 q724 q725
XSPLIT364 LSmitll_SPLIT 364 q726 q727
XSPLIT365 LSmitll_SPLIT 365 q728 q729
XSPLIT366 LSmitll_SPLIT 366 q730 q731
XSPLIT367 LSmitll_SPLIT 367 q732 q733
XSPLIT368 LSmitll_SPLIT 368 q734 q735
XSPLIT369 LSmitll_SPLIT 369 q736 q737
XSPLIT370 LSmitll_SPLIT 370 q738 q739
XSPLIT371 LSmitll_SPLIT 371 q740 q741
XSPLIT372 LSmitll_SPLIT 372 q742 q743
XSPLIT373 LSmitll_SPLIT 373 q744 q745
XSPLIT374 LSmitll_SPLIT 374 q746 q747
XSPLIT375 LSmitll_SPLIT 375 q748 q749
XSPLIT376 LSmitll_SPLIT 376 q750 q751
XSPLIT377 LSmitll_SPLIT 377 q752 q753
XSPLIT378 LSmitll_SPLIT 378 q754 q755
XSPLIT379 LSmitll_SPLIT 379 q756 q757
XSPLIT380 LSmitll_SPLIT 380 q758 q759
XSPLIT381 LSmitll_SPLIT 381 q760 q761
XSPLIT382 LSmitll_SPLIT 382 q762 q763
XSPLIT383 LSmitll_SPLIT 383 q764 q765
XSPLIT384 LSmitll_SPLIT 384 q766 q767
XSPLIT385 LSmitll_SPLIT 385 q768 q769
XSPLIT386 LSmitll_SPLIT 386 q770 q771
XSPLIT387 LSmitll_SPLIT 387 q772 q773
XSPLIT388 LSmitll_SPLIT 388 q774 q775
XSPLIT389 LSmitll_SPLIT 389 q776 q777
XSPLIT390 LSmitll_SPLIT 390 q778 q779
XSPLIT391 LSmitll_SPLIT 391 q780 q781
XSPLIT392 LSmitll_SPLIT 392 q782 q783
XSPLIT393 LSmitll_SPLIT 393 q784 q785
XSPLIT394 LSmitll_SPLIT 394 q786 q787
XSPLIT395 LSmitll_SPLIT 395 q788 q789
XSPLIT396 LSmitll_SPLIT 396 q790 q791
XSPLIT397 LSmitll_SPLIT 397 q792 q793
XSPLIT398 LSmitll_SPLIT 398 q794 q795
XSPLIT399 LSmitll_SPLIT 399 q796 q797
XSPLIT400 LSmitll_SPLIT 400 q798 q799
XSPLIT401 LSmitll_SPLIT 401 q800 q801
XSPLIT402 LSmitll_SPLIT 402 q802 q803
XSPLIT403 LSmitll_SPLIT 403 q804 q805
XSPLIT404 LSmitll_SPLIT 404 q806 q807
XSPLIT405 LSmitll_SPLIT 405 q808 q809
XSPLIT406 LSmitll_SPLIT 406 q810 q811
XSPLIT407 LSmitll_SPLIT 407 q812 q813
XSPLIT408 LSmitll_SPLIT 408 q814 q815
XSPLIT409 LSmitll_SPLIT 409 q816 q817
XSPLIT410 LSmitll_SPLIT 410 q818 q819
XSPLIT411 LSmitll_SPLIT 411 q820 q821
XSPLIT412 LSmitll_SPLIT 412 q822 q823
XSPLIT413 LSmitll_SPLIT 413 q824 q825
XSPLIT414 LSmitll_SPLIT 414 q826 q827
XSPLIT415 LSmitll_SPLIT 415 q828 q829
XSPLIT416 LSmitll_SPLIT 416 q830 q831
XSPLIT417 LSmitll_SPLIT 417 q832 q833
XSPLIT418 LSmitll_SPLIT 418 q834 q835
XSPLIT419 LSmitll_SPLIT 419 q836 q837
XSPLIT420 LSmitll_SPLIT 420 q838 q839
XSPLIT421 LSmitll_SPLIT 421 q840 q841
XSPLIT422 LSmitll_SPLIT 422 q842 q843
XSPLIT423 LSmitll_SPLIT 423 q844 q845
XSPLIT424 LSmitll_SPLIT 424 q846 q847
XSPLIT425 LSmitll_SPLIT 425 q848 q849
XSPLIT426 LSmitll_SPLIT 426 q850 q851
XSPLIT427 LSmitll_SPLIT 427 q852 q853
XSPLIT428 LSmitll_SPLIT 428 q854 q855
XSPLIT429 LSmitll_SPLIT 429 q856 q857
XSPLIT430 LSmitll_SPLIT 430 q858 q859
XSPLIT431 LSmitll_SPLIT 431 q860 q861
XSPLIT432 LSmitll_SPLIT 432 q862 q863
XSPLIT433 LSmitll_SPLIT 433 q864 q865
XSPLIT434 LSmitll_SPLIT 434 q866 q867
XSPLIT435 LSmitll_SPLIT 435 q868 q869
XSPLIT436 LSmitll_SPLIT 436 q870 q871
XSPLIT437 LSmitll_SPLIT 437 q872 q873
XSPLIT438 LSmitll_SPLIT 438 q874 q875
XSPLIT439 LSmitll_SPLIT 439 q876 q877
XSPLIT440 LSmitll_SPLIT 440 q878 q879
XSPLIT441 LSmitll_SPLIT 441 q880 q881
XSPLIT442 LSmitll_SPLIT 442 q882 q883
XSPLIT443 LSmitll_SPLIT 443 q884 q885
XSPLIT444 LSmitll_SPLIT 444 q886 q887
XSPLIT445 LSmitll_SPLIT 445 q888 q889
XSPLIT446 LSmitll_SPLIT 446 q890 q891
XSPLIT447 LSmitll_SPLIT 447 q892 q893
XSPLIT448 LSmitll_SPLIT 448 q894 q895
XSPLIT449 LSmitll_SPLIT 449 q896 q897
XSPLIT450 LSmitll_SPLIT 450 q898 q899
XSPLIT451 LSmitll_SPLIT 451 q900 q901
XSPLIT452 LSmitll_SPLIT 452 q902 q903
XSPLIT453 LSmitll_SPLIT 453 q904 q905
XSPLIT454 LSmitll_SPLIT 454 q906 q907
XSPLIT455 LSmitll_SPLIT 455 q908 q909
XSPLIT456 LSmitll_SPLIT 456 q910 q911
XSPLIT457 LSmitll_SPLIT 457 q912 q913
XSPLIT458 LSmitll_SPLIT 458 q914 q915
XSPLIT459 LSmitll_SPLIT 459 q916 q917
XSPLIT460 LSmitll_SPLIT 460 q918 q919
XSPLIT461 LSmitll_SPLIT 461 q920 q921
XSPLIT462 LSmitll_SPLIT 462 q922 q923
XSPLIT463 LSmitll_SPLIT 463 q924 q925
XSPLIT464 LSmitll_SPLIT 464 q926 q927
XSPLIT465 LSmitll_SPLIT 465 q928 q929
XSPLIT466 LSmitll_SPLIT 466 q930 q931
XSPLIT467 LSmitll_SPLIT 467 q932 q933
XSPLIT468 LSmitll_SPLIT 468 q934 q935
XSPLIT469 LSmitll_SPLIT 469 q936 q937
XSPLIT470 LSmitll_SPLIT 470 q938 q939
XSPLIT471 LSmitll_SPLIT 471 q940 q941
XSPLIT472 LSmitll_SPLIT 472 q942 q943
XSPLIT473 LSmitll_SPLIT 473 q944 q945
XSPLIT474 LSmitll_SPLIT 474 q946 q947
XSPLIT475 LSmitll_SPLIT 475 q948 q949
XSPLIT476 LSmitll_SPLIT 476 q950 q951
XSPLIT477 LSmitll_SPLIT 477 q952 q953
XSPLIT478 LSmitll_SPLIT 478 q954 q955
XSPLIT479 LSmitll_SPLIT 479 q956 q957
XSPLIT480 LSmitll_SPLIT 480 q958 q959
XSPLIT481 LSmitll_SPLIT 481 q960 q961
XSPLIT482 LSmitll_SPLIT 482 q962 q963
XSPLIT483 LSmitll_SPLIT 483 q964 q965
XSPLIT484 LSmitll_SPLIT 484 q966 q967
XSPLIT485 LSmitll_SPLIT 485 q968 q969
XSPLIT486 LSmitll_SPLIT 486 q970 q971
XSPLIT487 LSmitll_SPLIT 487 q972 q973
XSPLIT488 LSmitll_SPLIT 488 q974 q975
XSPLIT489 LSmitll_SPLIT 489 q976 q977
XSPLIT490 LSmitll_SPLIT 490 q978 q979
XSPLIT491 LSmitll_SPLIT 491 q980 q981
XSPLIT492 LSmitll_SPLIT 492 q982 q983
XSPLIT493 LSmitll_SPLIT 493 q984 q985
XSPLIT494 LSmitll_SPLIT 494 q986 q987
XSPLIT495 LSmitll_SPLIT 495 q988 q989
XSPLIT496 LSmitll_SPLIT 496 q990 q991
XSPLIT497 LSmitll_SPLIT 497 q992 q993
XSPLIT498 LSmitll_SPLIT 498 q994 q995
XSPLIT499 LSmitll_SPLIT 499 q996 q997
XSPLIT500 LSmitll_SPLIT 500 q998 q999
XSPLIT501 LSmitll_SPLIT 501 q1000 q1001
XSPLIT502 LSmitll_SPLIT 502 q1002 q1003
XSPLIT503 LSmitll_SPLIT 503 q1004 q1005
XSPLIT504 LSmitll_SPLIT 504 q1006 q1007
XSPLIT505 LSmitll_SPLIT 505 q1008 q1009
XSPLIT506 LSmitll_SPLIT 506 q1010 q1011
XSPLIT507 LSmitll_SPLIT 507 q1012 q1013
XSPLIT508 LSmitll_SPLIT 508 q1014 q1015
XSPLIT509 LSmitll_SPLIT 509 q1016 q1017
XSPLIT510 LSmitll_SPLIT 510 q1018 q1019
XSPLIT511 LSmitll_SPLIT 511 q1020 q1021
XSPLIT512 LSmitll_SPLIT 512 q1022 q1023
.ends 1_to_1024_split

.subckt 1_to_2048_split a q0 q1 q2 q3 q4 q5 q6 q7 q8 q9 q10 q11 q12 q13 q14 q15 q16 q17 q18 q19 q20 q21 q22 q23 q24 q25 q26 q27 q28 q29 q30 q31 q32 q33 q34 q35 q36 q37 q38 q39 q40 q41 q42 q43 q44 q45 q46 q47 q48 q49 q50 q51 q52 q53 q54 q55 q56 q57 q58 q59 q60 q61 q62 q63 q64 q65 q66 q67 q68 q69 q70 q71 q72 q73 q74 q75 q76 q77 q78 q79 q80 q81 q82 q83 q84 q85 q86 q87 q88 q89 q90 q91 q92 q93 q94 q95 q96 q97 q98 q99 q100 q101 q102 q103 q104 q105 q106 q107 q108 q109 q110 q111 q112 q113 q114 q115 q116 q117 q118 q119 q120 q121 q122 q123 q124 q125 q126 q127 q128 q129 q130 q131 q132 q133 q134 q135 q136 q137 q138 q139 q140 q141 q142 q143 q144 q145 q146 q147 q148 q149 q150 q151 q152 q153 q154 q155 q156 q157 q158 q159 q160 q161 q162 q163 q164 q165 q166 q167 q168 q169 q170 q171 q172 q173 q174 q175 q176 q177 q178 q179 q180 q181 q182 q183 q184 q185 q186 q187 q188 q189 q190 q191 q192 q193 q194 q195 q196 q197 q198 q199 q200 q201 q202 q203 q204 q205 q206 q207 q208 q209 q210 q211 q212 q213 q214 q215 q216 q217 q218 q219 q220 q221 q222 q223 q224 q225 q226 q227 q228 q229 q230 q231 q232 q233 q234 q235 q236 q237 q238 q239 q240 q241 q242 q243 q244 q245 q246 q247 q248 q249 q250 q251 q252 q253 q254 q255 q256 q257 q258 q259 q260 q261 q262 q263 q264 q265 q266 q267 q268 q269 q270 q271 q272 q273 q274 q275 q276 q277 q278 q279 q280 q281 q282 q283 q284 q285 q286 q287 q288 q289 q290 q291 q292 q293 q294 q295 q296 q297 q298 q299 q300 q301 q302 q303 q304 q305 q306 q307 q308 q309 q310 q311 q312 q313 q314 q315 q316 q317 q318 q319 q320 q321 q322 q323 q324 q325 q326 q327 q328 q329 q330 q331 q332 q333 q334 q335 q336 q337 q338 q339 q340 q341 q342 q343 q344 q345 q346 q347 q348 q349 q350 q351 q352 q353 q354 q355 q356 q357 q358 q359 q360 q361 q362 q363 q364 q365 q366 q367 q368 q369 q370 q371 q372 q373 q374 q375 q376 q377 q378 q379 q380 q381 q382 q383 q384 q385 q386 q387 q388 q389 q390 q391 q392 q393 q394 q395 q396 q397 q398 q399 q400 q401 q402 q403 q404 q405 q406 q407 q408 q409 q410 q411 q412 q413 q414 q415 q416 q417 q418 q419 q420 q421 q422 q423 q424 q425 q426 q427 q428 q429 q430 q431 q432 q433 q434 q435 q436 q437 q438 q439 q440 q441 q442 q443 q444 q445 q446 q447 q448 q449 q450 q451 q452 q453 q454 q455 q456 q457 q458 q459 q460 q461 q462 q463 q464 q465 q466 q467 q468 q469 q470 q471 q472 q473 q474 q475 q476 q477 q478 q479 q480 q481 q482 q483 q484 q485 q486 q487 q488 q489 q490 q491 q492 q493 q494 q495 q496 q497 q498 q499 q500 q501 q502 q503 q504 q505 q506 q507 q508 q509 q510 q511 q512 q513 q514 q515 q516 q517 q518 q519 q520 q521 q522 q523 q524 q525 q526 q527 q528 q529 q530 q531 q532 q533 q534 q535 q536 q537 q538 q539 q540 q541 q542 q543 q544 q545 q546 q547 q548 q549 q550 q551 q552 q553 q554 q555 q556 q557 q558 q559 q560 q561 q562 q563 q564 q565 q566 q567 q568 q569 q570 q571 q572 q573 q574 q575 q576 q577 q578 q579 q580 q581 q582 q583 q584 q585 q586 q587 q588 q589 q590 q591 q592 q593 q594 q595 q596 q597 q598 q599 q600 q601 q602 q603 q604 q605 q606 q607 q608 q609 q610 q611 q612 q613 q614 q615 q616 q617 q618 q619 q620 q621 q622 q623 q624 q625 q626 q627 q628 q629 q630 q631 q632 q633 q634 q635 q636 q637 q638 q639 q640 q641 q642 q643 q644 q645 q646 q647 q648 q649 q650 q651 q652 q653 q654 q655 q656 q657 q658 q659 q660 q661 q662 q663 q664 q665 q666 q667 q668 q669 q670 q671 q672 q673 q674 q675 q676 q677 q678 q679 q680 q681 q682 q683 q684 q685 q686 q687 q688 q689 q690 q691 q692 q693 q694 q695 q696 q697 q698 q699 q700 q701 q702 q703 q704 q705 q706 q707 q708 q709 q710 q711 q712 q713 q714 q715 q716 q717 q718 q719 q720 q721 q722 q723 q724 q725 q726 q727 q728 q729 q730 q731 q732 q733 q734 q735 q736 q737 q738 q739 q740 q741 q742 q743 q744 q745 q746 q747 q748 q749 q750 q751 q752 q753 q754 q755 q756 q757 q758 q759 q760 q761 q762 q763 q764 q765 q766 q767 q768 q769 q770 q771 q772 q773 q774 q775 q776 q777 q778 q779 q780 q781 q782 q783 q784 q785 q786 q787 q788 q789 q790 q791 q792 q793 q794 q795 q796 q797 q798 q799 q800 q801 q802 q803 q804 q805 q806 q807 q808 q809 q810 q811 q812 q813 q814 q815 q816 q817 q818 q819 q820 q821 q822 q823 q824 q825 q826 q827 q828 q829 q830 q831 q832 q833 q834 q835 q836 q837 q838 q839 q840 q841 q842 q843 q844 q845 q846 q847 q848 q849 q850 q851 q852 q853 q854 q855 q856 q857 q858 q859 q860 q861 q862 q863 q864 q865 q866 q867 q868 q869 q870 q871 q872 q873 q874 q875 q876 q877 q878 q879 q880 q881 q882 q883 q884 q885 q886 q887 q888 q889 q890 q891 q892 q893 q894 q895 q896 q897 q898 q899 q900 q901 q902 q903 q904 q905 q906 q907 q908 q909 q910 q911 q912 q913 q914 q915 q916 q917 q918 q919 q920 q921 q922 q923 q924 q925 q926 q927 q928 q929 q930 q931 q932 q933 q934 q935 q936 q937 q938 q939 q940 q941 q942 q943 q944 q945 q946 q947 q948 q949 q950 q951 q952 q953 q954 q955 q956 q957 q958 q959 q960 q961 q962 q963 q964 q965 q966 q967 q968 q969 q970 q971 q972 q973 q974 q975 q976 q977 q978 q979 q980 q981 q982 q983 q984 q985 q986 q987 q988 q989 q990 q991 q992 q993 q994 q995 q996 q997 q998 q999 q1000 q1001 q1002 q1003 q1004 q1005 q1006 q1007 q1008 q1009 q1010 q1011 q1012 q1013 q1014 q1015 q1016 q1017 q1018 q1019 q1020 q1021 q1022 q1023 q1024 q1025 q1026 q1027 q1028 q1029 q1030 q1031 q1032 q1033 q1034 q1035 q1036 q1037 q1038 q1039 q1040 q1041 q1042 q1043 q1044 q1045 q1046 q1047 q1048 q1049 q1050 q1051 q1052 q1053 q1054 q1055 q1056 q1057 q1058 q1059 q1060 q1061 q1062 q1063 q1064 q1065 q1066 q1067 q1068 q1069 q1070 q1071 q1072 q1073 q1074 q1075 q1076 q1077 q1078 q1079 q1080 q1081 q1082 q1083 q1084 q1085 q1086 q1087 q1088 q1089 q1090 q1091 q1092 q1093 q1094 q1095 q1096 q1097 q1098 q1099 q1100 q1101 q1102 q1103 q1104 q1105 q1106 q1107 q1108 q1109 q1110 q1111 q1112 q1113 q1114 q1115 q1116 q1117 q1118 q1119 q1120 q1121 q1122 q1123 q1124 q1125 q1126 q1127 q1128 q1129 q1130 q1131 q1132 q1133 q1134 q1135 q1136 q1137 q1138 q1139 q1140 q1141 q1142 q1143 q1144 q1145 q1146 q1147 q1148 q1149 q1150 q1151 q1152 q1153 q1154 q1155 q1156 q1157 q1158 q1159 q1160 q1161 q1162 q1163 q1164 q1165 q1166 q1167 q1168 q1169 q1170 q1171 q1172 q1173 q1174 q1175 q1176 q1177 q1178 q1179 q1180 q1181 q1182 q1183 q1184 q1185 q1186 q1187 q1188 q1189 q1190 q1191 q1192 q1193 q1194 q1195 q1196 q1197 q1198 q1199 q1200 q1201 q1202 q1203 q1204 q1205 q1206 q1207 q1208 q1209 q1210 q1211 q1212 q1213 q1214 q1215 q1216 q1217 q1218 q1219 q1220 q1221 q1222 q1223 q1224 q1225 q1226 q1227 q1228 q1229 q1230 q1231 q1232 q1233 q1234 q1235 q1236 q1237 q1238 q1239 q1240 q1241 q1242 q1243 q1244 q1245 q1246 q1247 q1248 q1249 q1250 q1251 q1252 q1253 q1254 q1255 q1256 q1257 q1258 q1259 q1260 q1261 q1262 q1263 q1264 q1265 q1266 q1267 q1268 q1269 q1270 q1271 q1272 q1273 q1274 q1275 q1276 q1277 q1278 q1279 q1280 q1281 q1282 q1283 q1284 q1285 q1286 q1287 q1288 q1289 q1290 q1291 q1292 q1293 q1294 q1295 q1296 q1297 q1298 q1299 q1300 q1301 q1302 q1303 q1304 q1305 q1306 q1307 q1308 q1309 q1310 q1311 q1312 q1313 q1314 q1315 q1316 q1317 q1318 q1319 q1320 q1321 q1322 q1323 q1324 q1325 q1326 q1327 q1328 q1329 q1330 q1331 q1332 q1333 q1334 q1335 q1336 q1337 q1338 q1339 q1340 q1341 q1342 q1343 q1344 q1345 q1346 q1347 q1348 q1349 q1350 q1351 q1352 q1353 q1354 q1355 q1356 q1357 q1358 q1359 q1360 q1361 q1362 q1363 q1364 q1365 q1366 q1367 q1368 q1369 q1370 q1371 q1372 q1373 q1374 q1375 q1376 q1377 q1378 q1379 q1380 q1381 q1382 q1383 q1384 q1385 q1386 q1387 q1388 q1389 q1390 q1391 q1392 q1393 q1394 q1395 q1396 q1397 q1398 q1399 q1400 q1401 q1402 q1403 q1404 q1405 q1406 q1407 q1408 q1409 q1410 q1411 q1412 q1413 q1414 q1415 q1416 q1417 q1418 q1419 q1420 q1421 q1422 q1423 q1424 q1425 q1426 q1427 q1428 q1429 q1430 q1431 q1432 q1433 q1434 q1435 q1436 q1437 q1438 q1439 q1440 q1441 q1442 q1443 q1444 q1445 q1446 q1447 q1448 q1449 q1450 q1451 q1452 q1453 q1454 q1455 q1456 q1457 q1458 q1459 q1460 q1461 q1462 q1463 q1464 q1465 q1466 q1467 q1468 q1469 q1470 q1471 q1472 q1473 q1474 q1475 q1476 q1477 q1478 q1479 q1480 q1481 q1482 q1483 q1484 q1485 q1486 q1487 q1488 q1489 q1490 q1491 q1492 q1493 q1494 q1495 q1496 q1497 q1498 q1499 q1500 q1501 q1502 q1503 q1504 q1505 q1506 q1507 q1508 q1509 q1510 q1511 q1512 q1513 q1514 q1515 q1516 q1517 q1518 q1519 q1520 q1521 q1522 q1523 q1524 q1525 q1526 q1527 q1528 q1529 q1530 q1531 q1532 q1533 q1534 q1535 q1536 q1537 q1538 q1539 q1540 q1541 q1542 q1543 q1544 q1545 q1546 q1547 q1548 q1549 q1550 q1551 q1552 q1553 q1554 q1555 q1556 q1557 q1558 q1559 q1560 q1561 q1562 q1563 q1564 q1565 q1566 q1567 q1568 q1569 q1570 q1571 q1572 q1573 q1574 q1575 q1576 q1577 q1578 q1579 q1580 q1581 q1582 q1583 q1584 q1585 q1586 q1587 q1588 q1589 q1590 q1591 q1592 q1593 q1594 q1595 q1596 q1597 q1598 q1599 q1600 q1601 q1602 q1603 q1604 q1605 q1606 q1607 q1608 q1609 q1610 q1611 q1612 q1613 q1614 q1615 q1616 q1617 q1618 q1619 q1620 q1621 q1622 q1623 q1624 q1625 q1626 q1627 q1628 q1629 q1630 q1631 q1632 q1633 q1634 q1635 q1636 q1637 q1638 q1639 q1640 q1641 q1642 q1643 q1644 q1645 q1646 q1647 q1648 q1649 q1650 q1651 q1652 q1653 q1654 q1655 q1656 q1657 q1658 q1659 q1660 q1661 q1662 q1663 q1664 q1665 q1666 q1667 q1668 q1669 q1670 q1671 q1672 q1673 q1674 q1675 q1676 q1677 q1678 q1679 q1680 q1681 q1682 q1683 q1684 q1685 q1686 q1687 q1688 q1689 q1690 q1691 q1692 q1693 q1694 q1695 q1696 q1697 q1698 q1699 q1700 q1701 q1702 q1703 q1704 q1705 q1706 q1707 q1708 q1709 q1710 q1711 q1712 q1713 q1714 q1715 q1716 q1717 q1718 q1719 q1720 q1721 q1722 q1723 q1724 q1725 q1726 q1727 q1728 q1729 q1730 q1731 q1732 q1733 q1734 q1735 q1736 q1737 q1738 q1739 q1740 q1741 q1742 q1743 q1744 q1745 q1746 q1747 q1748 q1749 q1750 q1751 q1752 q1753 q1754 q1755 q1756 q1757 q1758 q1759 q1760 q1761 q1762 q1763 q1764 q1765 q1766 q1767 q1768 q1769 q1770 q1771 q1772 q1773 q1774 q1775 q1776 q1777 q1778 q1779 q1780 q1781 q1782 q1783 q1784 q1785 q1786 q1787 q1788 q1789 q1790 q1791 q1792 q1793 q1794 q1795 q1796 q1797 q1798 q1799 q1800 q1801 q1802 q1803 q1804 q1805 q1806 q1807 q1808 q1809 q1810 q1811 q1812 q1813 q1814 q1815 q1816 q1817 q1818 q1819 q1820 q1821 q1822 q1823 q1824 q1825 q1826 q1827 q1828 q1829 q1830 q1831 q1832 q1833 q1834 q1835 q1836 q1837 q1838 q1839 q1840 q1841 q1842 q1843 q1844 q1845 q1846 q1847 q1848 q1849 q1850 q1851 q1852 q1853 q1854 q1855 q1856 q1857 q1858 q1859 q1860 q1861 q1862 q1863 q1864 q1865 q1866 q1867 q1868 q1869 q1870 q1871 q1872 q1873 q1874 q1875 q1876 q1877 q1878 q1879 q1880 q1881 q1882 q1883 q1884 q1885 q1886 q1887 q1888 q1889 q1890 q1891 q1892 q1893 q1894 q1895 q1896 q1897 q1898 q1899 q1900 q1901 q1902 q1903 q1904 q1905 q1906 q1907 q1908 q1909 q1910 q1911 q1912 q1913 q1914 q1915 q1916 q1917 q1918 q1919 q1920 q1921 q1922 q1923 q1924 q1925 q1926 q1927 q1928 q1929 q1930 q1931 q1932 q1933 q1934 q1935 q1936 q1937 q1938 q1939 q1940 q1941 q1942 q1943 q1944 q1945 q1946 q1947 q1948 q1949 q1950 q1951 q1952 q1953 q1954 q1955 q1956 q1957 q1958 q1959 q1960 q1961 q1962 q1963 q1964 q1965 q1966 q1967 q1968 q1969 q1970 q1971 q1972 q1973 q1974 q1975 q1976 q1977 q1978 q1979 q1980 q1981 q1982 q1983 q1984 q1985 q1986 q1987 q1988 q1989 q1990 q1991 q1992 q1993 q1994 q1995 q1996 q1997 q1998 q1999 q2000 q2001 q2002 q2003 q2004 q2005 q2006 q2007 q2008 q2009 q2010 q2011 q2012 q2013 q2014 q2015 q2016 q2017 q2018 q2019 q2020 q2021 q2022 q2023 q2024 q2025 q2026 q2027 q2028 q2029 q2030 q2031 q2032 q2033 q2034 q2035 q2036 q2037 q2038 q2039 q2040 q2041 q2042 q2043 q2044 q2045 q2046 q2047 
XSPLIT_1024 1_to_1024_split a 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921 922 923 924 925 926 927 928 929 930 931 932 933 934 935 936 937 938 939 940 941 942 943 944 945 946 947 948 949 950 951 952 953 954 955 956 957 958 959 960 961 962 963 964 965 966 967 968 969 970 971 972 973 974 975 976 977 978 979 980 981 982 983 984 985 986 987 988 989 990 991 992 993 994 995 996 997 998 999 1000 1001 1002 1003 1004 1005 1006 1007 1008 1009 1010 1011 1012 1013 1014 1015 1016 1017 1018 1019 1020 1021 1022 1023 1024 
XSPLIT1 LSmitll_SPLIT 1 q0 q1
XSPLIT2 LSmitll_SPLIT 2 q2 q3
XSPLIT3 LSmitll_SPLIT 3 q4 q5
XSPLIT4 LSmitll_SPLIT 4 q6 q7
XSPLIT5 LSmitll_SPLIT 5 q8 q9
XSPLIT6 LSmitll_SPLIT 6 q10 q11
XSPLIT7 LSmitll_SPLIT 7 q12 q13
XSPLIT8 LSmitll_SPLIT 8 q14 q15
XSPLIT9 LSmitll_SPLIT 9 q16 q17
XSPLIT10 LSmitll_SPLIT 10 q18 q19
XSPLIT11 LSmitll_SPLIT 11 q20 q21
XSPLIT12 LSmitll_SPLIT 12 q22 q23
XSPLIT13 LSmitll_SPLIT 13 q24 q25
XSPLIT14 LSmitll_SPLIT 14 q26 q27
XSPLIT15 LSmitll_SPLIT 15 q28 q29
XSPLIT16 LSmitll_SPLIT 16 q30 q31
XSPLIT17 LSmitll_SPLIT 17 q32 q33
XSPLIT18 LSmitll_SPLIT 18 q34 q35
XSPLIT19 LSmitll_SPLIT 19 q36 q37
XSPLIT20 LSmitll_SPLIT 20 q38 q39
XSPLIT21 LSmitll_SPLIT 21 q40 q41
XSPLIT22 LSmitll_SPLIT 22 q42 q43
XSPLIT23 LSmitll_SPLIT 23 q44 q45
XSPLIT24 LSmitll_SPLIT 24 q46 q47
XSPLIT25 LSmitll_SPLIT 25 q48 q49
XSPLIT26 LSmitll_SPLIT 26 q50 q51
XSPLIT27 LSmitll_SPLIT 27 q52 q53
XSPLIT28 LSmitll_SPLIT 28 q54 q55
XSPLIT29 LSmitll_SPLIT 29 q56 q57
XSPLIT30 LSmitll_SPLIT 30 q58 q59
XSPLIT31 LSmitll_SPLIT 31 q60 q61
XSPLIT32 LSmitll_SPLIT 32 q62 q63
XSPLIT33 LSmitll_SPLIT 33 q64 q65
XSPLIT34 LSmitll_SPLIT 34 q66 q67
XSPLIT35 LSmitll_SPLIT 35 q68 q69
XSPLIT36 LSmitll_SPLIT 36 q70 q71
XSPLIT37 LSmitll_SPLIT 37 q72 q73
XSPLIT38 LSmitll_SPLIT 38 q74 q75
XSPLIT39 LSmitll_SPLIT 39 q76 q77
XSPLIT40 LSmitll_SPLIT 40 q78 q79
XSPLIT41 LSmitll_SPLIT 41 q80 q81
XSPLIT42 LSmitll_SPLIT 42 q82 q83
XSPLIT43 LSmitll_SPLIT 43 q84 q85
XSPLIT44 LSmitll_SPLIT 44 q86 q87
XSPLIT45 LSmitll_SPLIT 45 q88 q89
XSPLIT46 LSmitll_SPLIT 46 q90 q91
XSPLIT47 LSmitll_SPLIT 47 q92 q93
XSPLIT48 LSmitll_SPLIT 48 q94 q95
XSPLIT49 LSmitll_SPLIT 49 q96 q97
XSPLIT50 LSmitll_SPLIT 50 q98 q99
XSPLIT51 LSmitll_SPLIT 51 q100 q101
XSPLIT52 LSmitll_SPLIT 52 q102 q103
XSPLIT53 LSmitll_SPLIT 53 q104 q105
XSPLIT54 LSmitll_SPLIT 54 q106 q107
XSPLIT55 LSmitll_SPLIT 55 q108 q109
XSPLIT56 LSmitll_SPLIT 56 q110 q111
XSPLIT57 LSmitll_SPLIT 57 q112 q113
XSPLIT58 LSmitll_SPLIT 58 q114 q115
XSPLIT59 LSmitll_SPLIT 59 q116 q117
XSPLIT60 LSmitll_SPLIT 60 q118 q119
XSPLIT61 LSmitll_SPLIT 61 q120 q121
XSPLIT62 LSmitll_SPLIT 62 q122 q123
XSPLIT63 LSmitll_SPLIT 63 q124 q125
XSPLIT64 LSmitll_SPLIT 64 q126 q127
XSPLIT65 LSmitll_SPLIT 65 q128 q129
XSPLIT66 LSmitll_SPLIT 66 q130 q131
XSPLIT67 LSmitll_SPLIT 67 q132 q133
XSPLIT68 LSmitll_SPLIT 68 q134 q135
XSPLIT69 LSmitll_SPLIT 69 q136 q137
XSPLIT70 LSmitll_SPLIT 70 q138 q139
XSPLIT71 LSmitll_SPLIT 71 q140 q141
XSPLIT72 LSmitll_SPLIT 72 q142 q143
XSPLIT73 LSmitll_SPLIT 73 q144 q145
XSPLIT74 LSmitll_SPLIT 74 q146 q147
XSPLIT75 LSmitll_SPLIT 75 q148 q149
XSPLIT76 LSmitll_SPLIT 76 q150 q151
XSPLIT77 LSmitll_SPLIT 77 q152 q153
XSPLIT78 LSmitll_SPLIT 78 q154 q155
XSPLIT79 LSmitll_SPLIT 79 q156 q157
XSPLIT80 LSmitll_SPLIT 80 q158 q159
XSPLIT81 LSmitll_SPLIT 81 q160 q161
XSPLIT82 LSmitll_SPLIT 82 q162 q163
XSPLIT83 LSmitll_SPLIT 83 q164 q165
XSPLIT84 LSmitll_SPLIT 84 q166 q167
XSPLIT85 LSmitll_SPLIT 85 q168 q169
XSPLIT86 LSmitll_SPLIT 86 q170 q171
XSPLIT87 LSmitll_SPLIT 87 q172 q173
XSPLIT88 LSmitll_SPLIT 88 q174 q175
XSPLIT89 LSmitll_SPLIT 89 q176 q177
XSPLIT90 LSmitll_SPLIT 90 q178 q179
XSPLIT91 LSmitll_SPLIT 91 q180 q181
XSPLIT92 LSmitll_SPLIT 92 q182 q183
XSPLIT93 LSmitll_SPLIT 93 q184 q185
XSPLIT94 LSmitll_SPLIT 94 q186 q187
XSPLIT95 LSmitll_SPLIT 95 q188 q189
XSPLIT96 LSmitll_SPLIT 96 q190 q191
XSPLIT97 LSmitll_SPLIT 97 q192 q193
XSPLIT98 LSmitll_SPLIT 98 q194 q195
XSPLIT99 LSmitll_SPLIT 99 q196 q197
XSPLIT100 LSmitll_SPLIT 100 q198 q199
XSPLIT101 LSmitll_SPLIT 101 q200 q201
XSPLIT102 LSmitll_SPLIT 102 q202 q203
XSPLIT103 LSmitll_SPLIT 103 q204 q205
XSPLIT104 LSmitll_SPLIT 104 q206 q207
XSPLIT105 LSmitll_SPLIT 105 q208 q209
XSPLIT106 LSmitll_SPLIT 106 q210 q211
XSPLIT107 LSmitll_SPLIT 107 q212 q213
XSPLIT108 LSmitll_SPLIT 108 q214 q215
XSPLIT109 LSmitll_SPLIT 109 q216 q217
XSPLIT110 LSmitll_SPLIT 110 q218 q219
XSPLIT111 LSmitll_SPLIT 111 q220 q221
XSPLIT112 LSmitll_SPLIT 112 q222 q223
XSPLIT113 LSmitll_SPLIT 113 q224 q225
XSPLIT114 LSmitll_SPLIT 114 q226 q227
XSPLIT115 LSmitll_SPLIT 115 q228 q229
XSPLIT116 LSmitll_SPLIT 116 q230 q231
XSPLIT117 LSmitll_SPLIT 117 q232 q233
XSPLIT118 LSmitll_SPLIT 118 q234 q235
XSPLIT119 LSmitll_SPLIT 119 q236 q237
XSPLIT120 LSmitll_SPLIT 120 q238 q239
XSPLIT121 LSmitll_SPLIT 121 q240 q241
XSPLIT122 LSmitll_SPLIT 122 q242 q243
XSPLIT123 LSmitll_SPLIT 123 q244 q245
XSPLIT124 LSmitll_SPLIT 124 q246 q247
XSPLIT125 LSmitll_SPLIT 125 q248 q249
XSPLIT126 LSmitll_SPLIT 126 q250 q251
XSPLIT127 LSmitll_SPLIT 127 q252 q253
XSPLIT128 LSmitll_SPLIT 128 q254 q255
XSPLIT129 LSmitll_SPLIT 129 q256 q257
XSPLIT130 LSmitll_SPLIT 130 q258 q259
XSPLIT131 LSmitll_SPLIT 131 q260 q261
XSPLIT132 LSmitll_SPLIT 132 q262 q263
XSPLIT133 LSmitll_SPLIT 133 q264 q265
XSPLIT134 LSmitll_SPLIT 134 q266 q267
XSPLIT135 LSmitll_SPLIT 135 q268 q269
XSPLIT136 LSmitll_SPLIT 136 q270 q271
XSPLIT137 LSmitll_SPLIT 137 q272 q273
XSPLIT138 LSmitll_SPLIT 138 q274 q275
XSPLIT139 LSmitll_SPLIT 139 q276 q277
XSPLIT140 LSmitll_SPLIT 140 q278 q279
XSPLIT141 LSmitll_SPLIT 141 q280 q281
XSPLIT142 LSmitll_SPLIT 142 q282 q283
XSPLIT143 LSmitll_SPLIT 143 q284 q285
XSPLIT144 LSmitll_SPLIT 144 q286 q287
XSPLIT145 LSmitll_SPLIT 145 q288 q289
XSPLIT146 LSmitll_SPLIT 146 q290 q291
XSPLIT147 LSmitll_SPLIT 147 q292 q293
XSPLIT148 LSmitll_SPLIT 148 q294 q295
XSPLIT149 LSmitll_SPLIT 149 q296 q297
XSPLIT150 LSmitll_SPLIT 150 q298 q299
XSPLIT151 LSmitll_SPLIT 151 q300 q301
XSPLIT152 LSmitll_SPLIT 152 q302 q303
XSPLIT153 LSmitll_SPLIT 153 q304 q305
XSPLIT154 LSmitll_SPLIT 154 q306 q307
XSPLIT155 LSmitll_SPLIT 155 q308 q309
XSPLIT156 LSmitll_SPLIT 156 q310 q311
XSPLIT157 LSmitll_SPLIT 157 q312 q313
XSPLIT158 LSmitll_SPLIT 158 q314 q315
XSPLIT159 LSmitll_SPLIT 159 q316 q317
XSPLIT160 LSmitll_SPLIT 160 q318 q319
XSPLIT161 LSmitll_SPLIT 161 q320 q321
XSPLIT162 LSmitll_SPLIT 162 q322 q323
XSPLIT163 LSmitll_SPLIT 163 q324 q325
XSPLIT164 LSmitll_SPLIT 164 q326 q327
XSPLIT165 LSmitll_SPLIT 165 q328 q329
XSPLIT166 LSmitll_SPLIT 166 q330 q331
XSPLIT167 LSmitll_SPLIT 167 q332 q333
XSPLIT168 LSmitll_SPLIT 168 q334 q335
XSPLIT169 LSmitll_SPLIT 169 q336 q337
XSPLIT170 LSmitll_SPLIT 170 q338 q339
XSPLIT171 LSmitll_SPLIT 171 q340 q341
XSPLIT172 LSmitll_SPLIT 172 q342 q343
XSPLIT173 LSmitll_SPLIT 173 q344 q345
XSPLIT174 LSmitll_SPLIT 174 q346 q347
XSPLIT175 LSmitll_SPLIT 175 q348 q349
XSPLIT176 LSmitll_SPLIT 176 q350 q351
XSPLIT177 LSmitll_SPLIT 177 q352 q353
XSPLIT178 LSmitll_SPLIT 178 q354 q355
XSPLIT179 LSmitll_SPLIT 179 q356 q357
XSPLIT180 LSmitll_SPLIT 180 q358 q359
XSPLIT181 LSmitll_SPLIT 181 q360 q361
XSPLIT182 LSmitll_SPLIT 182 q362 q363
XSPLIT183 LSmitll_SPLIT 183 q364 q365
XSPLIT184 LSmitll_SPLIT 184 q366 q367
XSPLIT185 LSmitll_SPLIT 185 q368 q369
XSPLIT186 LSmitll_SPLIT 186 q370 q371
XSPLIT187 LSmitll_SPLIT 187 q372 q373
XSPLIT188 LSmitll_SPLIT 188 q374 q375
XSPLIT189 LSmitll_SPLIT 189 q376 q377
XSPLIT190 LSmitll_SPLIT 190 q378 q379
XSPLIT191 LSmitll_SPLIT 191 q380 q381
XSPLIT192 LSmitll_SPLIT 192 q382 q383
XSPLIT193 LSmitll_SPLIT 193 q384 q385
XSPLIT194 LSmitll_SPLIT 194 q386 q387
XSPLIT195 LSmitll_SPLIT 195 q388 q389
XSPLIT196 LSmitll_SPLIT 196 q390 q391
XSPLIT197 LSmitll_SPLIT 197 q392 q393
XSPLIT198 LSmitll_SPLIT 198 q394 q395
XSPLIT199 LSmitll_SPLIT 199 q396 q397
XSPLIT200 LSmitll_SPLIT 200 q398 q399
XSPLIT201 LSmitll_SPLIT 201 q400 q401
XSPLIT202 LSmitll_SPLIT 202 q402 q403
XSPLIT203 LSmitll_SPLIT 203 q404 q405
XSPLIT204 LSmitll_SPLIT 204 q406 q407
XSPLIT205 LSmitll_SPLIT 205 q408 q409
XSPLIT206 LSmitll_SPLIT 206 q410 q411
XSPLIT207 LSmitll_SPLIT 207 q412 q413
XSPLIT208 LSmitll_SPLIT 208 q414 q415
XSPLIT209 LSmitll_SPLIT 209 q416 q417
XSPLIT210 LSmitll_SPLIT 210 q418 q419
XSPLIT211 LSmitll_SPLIT 211 q420 q421
XSPLIT212 LSmitll_SPLIT 212 q422 q423
XSPLIT213 LSmitll_SPLIT 213 q424 q425
XSPLIT214 LSmitll_SPLIT 214 q426 q427
XSPLIT215 LSmitll_SPLIT 215 q428 q429
XSPLIT216 LSmitll_SPLIT 216 q430 q431
XSPLIT217 LSmitll_SPLIT 217 q432 q433
XSPLIT218 LSmitll_SPLIT 218 q434 q435
XSPLIT219 LSmitll_SPLIT 219 q436 q437
XSPLIT220 LSmitll_SPLIT 220 q438 q439
XSPLIT221 LSmitll_SPLIT 221 q440 q441
XSPLIT222 LSmitll_SPLIT 222 q442 q443
XSPLIT223 LSmitll_SPLIT 223 q444 q445
XSPLIT224 LSmitll_SPLIT 224 q446 q447
XSPLIT225 LSmitll_SPLIT 225 q448 q449
XSPLIT226 LSmitll_SPLIT 226 q450 q451
XSPLIT227 LSmitll_SPLIT 227 q452 q453
XSPLIT228 LSmitll_SPLIT 228 q454 q455
XSPLIT229 LSmitll_SPLIT 229 q456 q457
XSPLIT230 LSmitll_SPLIT 230 q458 q459
XSPLIT231 LSmitll_SPLIT 231 q460 q461
XSPLIT232 LSmitll_SPLIT 232 q462 q463
XSPLIT233 LSmitll_SPLIT 233 q464 q465
XSPLIT234 LSmitll_SPLIT 234 q466 q467
XSPLIT235 LSmitll_SPLIT 235 q468 q469
XSPLIT236 LSmitll_SPLIT 236 q470 q471
XSPLIT237 LSmitll_SPLIT 237 q472 q473
XSPLIT238 LSmitll_SPLIT 238 q474 q475
XSPLIT239 LSmitll_SPLIT 239 q476 q477
XSPLIT240 LSmitll_SPLIT 240 q478 q479
XSPLIT241 LSmitll_SPLIT 241 q480 q481
XSPLIT242 LSmitll_SPLIT 242 q482 q483
XSPLIT243 LSmitll_SPLIT 243 q484 q485
XSPLIT244 LSmitll_SPLIT 244 q486 q487
XSPLIT245 LSmitll_SPLIT 245 q488 q489
XSPLIT246 LSmitll_SPLIT 246 q490 q491
XSPLIT247 LSmitll_SPLIT 247 q492 q493
XSPLIT248 LSmitll_SPLIT 248 q494 q495
XSPLIT249 LSmitll_SPLIT 249 q496 q497
XSPLIT250 LSmitll_SPLIT 250 q498 q499
XSPLIT251 LSmitll_SPLIT 251 q500 q501
XSPLIT252 LSmitll_SPLIT 252 q502 q503
XSPLIT253 LSmitll_SPLIT 253 q504 q505
XSPLIT254 LSmitll_SPLIT 254 q506 q507
XSPLIT255 LSmitll_SPLIT 255 q508 q509
XSPLIT256 LSmitll_SPLIT 256 q510 q511
XSPLIT257 LSmitll_SPLIT 257 q512 q513
XSPLIT258 LSmitll_SPLIT 258 q514 q515
XSPLIT259 LSmitll_SPLIT 259 q516 q517
XSPLIT260 LSmitll_SPLIT 260 q518 q519
XSPLIT261 LSmitll_SPLIT 261 q520 q521
XSPLIT262 LSmitll_SPLIT 262 q522 q523
XSPLIT263 LSmitll_SPLIT 263 q524 q525
XSPLIT264 LSmitll_SPLIT 264 q526 q527
XSPLIT265 LSmitll_SPLIT 265 q528 q529
XSPLIT266 LSmitll_SPLIT 266 q530 q531
XSPLIT267 LSmitll_SPLIT 267 q532 q533
XSPLIT268 LSmitll_SPLIT 268 q534 q535
XSPLIT269 LSmitll_SPLIT 269 q536 q537
XSPLIT270 LSmitll_SPLIT 270 q538 q539
XSPLIT271 LSmitll_SPLIT 271 q540 q541
XSPLIT272 LSmitll_SPLIT 272 q542 q543
XSPLIT273 LSmitll_SPLIT 273 q544 q545
XSPLIT274 LSmitll_SPLIT 274 q546 q547
XSPLIT275 LSmitll_SPLIT 275 q548 q549
XSPLIT276 LSmitll_SPLIT 276 q550 q551
XSPLIT277 LSmitll_SPLIT 277 q552 q553
XSPLIT278 LSmitll_SPLIT 278 q554 q555
XSPLIT279 LSmitll_SPLIT 279 q556 q557
XSPLIT280 LSmitll_SPLIT 280 q558 q559
XSPLIT281 LSmitll_SPLIT 281 q560 q561
XSPLIT282 LSmitll_SPLIT 282 q562 q563
XSPLIT283 LSmitll_SPLIT 283 q564 q565
XSPLIT284 LSmitll_SPLIT 284 q566 q567
XSPLIT285 LSmitll_SPLIT 285 q568 q569
XSPLIT286 LSmitll_SPLIT 286 q570 q571
XSPLIT287 LSmitll_SPLIT 287 q572 q573
XSPLIT288 LSmitll_SPLIT 288 q574 q575
XSPLIT289 LSmitll_SPLIT 289 q576 q577
XSPLIT290 LSmitll_SPLIT 290 q578 q579
XSPLIT291 LSmitll_SPLIT 291 q580 q581
XSPLIT292 LSmitll_SPLIT 292 q582 q583
XSPLIT293 LSmitll_SPLIT 293 q584 q585
XSPLIT294 LSmitll_SPLIT 294 q586 q587
XSPLIT295 LSmitll_SPLIT 295 q588 q589
XSPLIT296 LSmitll_SPLIT 296 q590 q591
XSPLIT297 LSmitll_SPLIT 297 q592 q593
XSPLIT298 LSmitll_SPLIT 298 q594 q595
XSPLIT299 LSmitll_SPLIT 299 q596 q597
XSPLIT300 LSmitll_SPLIT 300 q598 q599
XSPLIT301 LSmitll_SPLIT 301 q600 q601
XSPLIT302 LSmitll_SPLIT 302 q602 q603
XSPLIT303 LSmitll_SPLIT 303 q604 q605
XSPLIT304 LSmitll_SPLIT 304 q606 q607
XSPLIT305 LSmitll_SPLIT 305 q608 q609
XSPLIT306 LSmitll_SPLIT 306 q610 q611
XSPLIT307 LSmitll_SPLIT 307 q612 q613
XSPLIT308 LSmitll_SPLIT 308 q614 q615
XSPLIT309 LSmitll_SPLIT 309 q616 q617
XSPLIT310 LSmitll_SPLIT 310 q618 q619
XSPLIT311 LSmitll_SPLIT 311 q620 q621
XSPLIT312 LSmitll_SPLIT 312 q622 q623
XSPLIT313 LSmitll_SPLIT 313 q624 q625
XSPLIT314 LSmitll_SPLIT 314 q626 q627
XSPLIT315 LSmitll_SPLIT 315 q628 q629
XSPLIT316 LSmitll_SPLIT 316 q630 q631
XSPLIT317 LSmitll_SPLIT 317 q632 q633
XSPLIT318 LSmitll_SPLIT 318 q634 q635
XSPLIT319 LSmitll_SPLIT 319 q636 q637
XSPLIT320 LSmitll_SPLIT 320 q638 q639
XSPLIT321 LSmitll_SPLIT 321 q640 q641
XSPLIT322 LSmitll_SPLIT 322 q642 q643
XSPLIT323 LSmitll_SPLIT 323 q644 q645
XSPLIT324 LSmitll_SPLIT 324 q646 q647
XSPLIT325 LSmitll_SPLIT 325 q648 q649
XSPLIT326 LSmitll_SPLIT 326 q650 q651
XSPLIT327 LSmitll_SPLIT 327 q652 q653
XSPLIT328 LSmitll_SPLIT 328 q654 q655
XSPLIT329 LSmitll_SPLIT 329 q656 q657
XSPLIT330 LSmitll_SPLIT 330 q658 q659
XSPLIT331 LSmitll_SPLIT 331 q660 q661
XSPLIT332 LSmitll_SPLIT 332 q662 q663
XSPLIT333 LSmitll_SPLIT 333 q664 q665
XSPLIT334 LSmitll_SPLIT 334 q666 q667
XSPLIT335 LSmitll_SPLIT 335 q668 q669
XSPLIT336 LSmitll_SPLIT 336 q670 q671
XSPLIT337 LSmitll_SPLIT 337 q672 q673
XSPLIT338 LSmitll_SPLIT 338 q674 q675
XSPLIT339 LSmitll_SPLIT 339 q676 q677
XSPLIT340 LSmitll_SPLIT 340 q678 q679
XSPLIT341 LSmitll_SPLIT 341 q680 q681
XSPLIT342 LSmitll_SPLIT 342 q682 q683
XSPLIT343 LSmitll_SPLIT 343 q684 q685
XSPLIT344 LSmitll_SPLIT 344 q686 q687
XSPLIT345 LSmitll_SPLIT 345 q688 q689
XSPLIT346 LSmitll_SPLIT 346 q690 q691
XSPLIT347 LSmitll_SPLIT 347 q692 q693
XSPLIT348 LSmitll_SPLIT 348 q694 q695
XSPLIT349 LSmitll_SPLIT 349 q696 q697
XSPLIT350 LSmitll_SPLIT 350 q698 q699
XSPLIT351 LSmitll_SPLIT 351 q700 q701
XSPLIT352 LSmitll_SPLIT 352 q702 q703
XSPLIT353 LSmitll_SPLIT 353 q704 q705
XSPLIT354 LSmitll_SPLIT 354 q706 q707
XSPLIT355 LSmitll_SPLIT 355 q708 q709
XSPLIT356 LSmitll_SPLIT 356 q710 q711
XSPLIT357 LSmitll_SPLIT 357 q712 q713
XSPLIT358 LSmitll_SPLIT 358 q714 q715
XSPLIT359 LSmitll_SPLIT 359 q716 q717
XSPLIT360 LSmitll_SPLIT 360 q718 q719
XSPLIT361 LSmitll_SPLIT 361 q720 q721
XSPLIT362 LSmitll_SPLIT 362 q722 q723
XSPLIT363 LSmitll_SPLIT 363 q724 q725
XSPLIT364 LSmitll_SPLIT 364 q726 q727
XSPLIT365 LSmitll_SPLIT 365 q728 q729
XSPLIT366 LSmitll_SPLIT 366 q730 q731
XSPLIT367 LSmitll_SPLIT 367 q732 q733
XSPLIT368 LSmitll_SPLIT 368 q734 q735
XSPLIT369 LSmitll_SPLIT 369 q736 q737
XSPLIT370 LSmitll_SPLIT 370 q738 q739
XSPLIT371 LSmitll_SPLIT 371 q740 q741
XSPLIT372 LSmitll_SPLIT 372 q742 q743
XSPLIT373 LSmitll_SPLIT 373 q744 q745
XSPLIT374 LSmitll_SPLIT 374 q746 q747
XSPLIT375 LSmitll_SPLIT 375 q748 q749
XSPLIT376 LSmitll_SPLIT 376 q750 q751
XSPLIT377 LSmitll_SPLIT 377 q752 q753
XSPLIT378 LSmitll_SPLIT 378 q754 q755
XSPLIT379 LSmitll_SPLIT 379 q756 q757
XSPLIT380 LSmitll_SPLIT 380 q758 q759
XSPLIT381 LSmitll_SPLIT 381 q760 q761
XSPLIT382 LSmitll_SPLIT 382 q762 q763
XSPLIT383 LSmitll_SPLIT 383 q764 q765
XSPLIT384 LSmitll_SPLIT 384 q766 q767
XSPLIT385 LSmitll_SPLIT 385 q768 q769
XSPLIT386 LSmitll_SPLIT 386 q770 q771
XSPLIT387 LSmitll_SPLIT 387 q772 q773
XSPLIT388 LSmitll_SPLIT 388 q774 q775
XSPLIT389 LSmitll_SPLIT 389 q776 q777
XSPLIT390 LSmitll_SPLIT 390 q778 q779
XSPLIT391 LSmitll_SPLIT 391 q780 q781
XSPLIT392 LSmitll_SPLIT 392 q782 q783
XSPLIT393 LSmitll_SPLIT 393 q784 q785
XSPLIT394 LSmitll_SPLIT 394 q786 q787
XSPLIT395 LSmitll_SPLIT 395 q788 q789
XSPLIT396 LSmitll_SPLIT 396 q790 q791
XSPLIT397 LSmitll_SPLIT 397 q792 q793
XSPLIT398 LSmitll_SPLIT 398 q794 q795
XSPLIT399 LSmitll_SPLIT 399 q796 q797
XSPLIT400 LSmitll_SPLIT 400 q798 q799
XSPLIT401 LSmitll_SPLIT 401 q800 q801
XSPLIT402 LSmitll_SPLIT 402 q802 q803
XSPLIT403 LSmitll_SPLIT 403 q804 q805
XSPLIT404 LSmitll_SPLIT 404 q806 q807
XSPLIT405 LSmitll_SPLIT 405 q808 q809
XSPLIT406 LSmitll_SPLIT 406 q810 q811
XSPLIT407 LSmitll_SPLIT 407 q812 q813
XSPLIT408 LSmitll_SPLIT 408 q814 q815
XSPLIT409 LSmitll_SPLIT 409 q816 q817
XSPLIT410 LSmitll_SPLIT 410 q818 q819
XSPLIT411 LSmitll_SPLIT 411 q820 q821
XSPLIT412 LSmitll_SPLIT 412 q822 q823
XSPLIT413 LSmitll_SPLIT 413 q824 q825
XSPLIT414 LSmitll_SPLIT 414 q826 q827
XSPLIT415 LSmitll_SPLIT 415 q828 q829
XSPLIT416 LSmitll_SPLIT 416 q830 q831
XSPLIT417 LSmitll_SPLIT 417 q832 q833
XSPLIT418 LSmitll_SPLIT 418 q834 q835
XSPLIT419 LSmitll_SPLIT 419 q836 q837
XSPLIT420 LSmitll_SPLIT 420 q838 q839
XSPLIT421 LSmitll_SPLIT 421 q840 q841
XSPLIT422 LSmitll_SPLIT 422 q842 q843
XSPLIT423 LSmitll_SPLIT 423 q844 q845
XSPLIT424 LSmitll_SPLIT 424 q846 q847
XSPLIT425 LSmitll_SPLIT 425 q848 q849
XSPLIT426 LSmitll_SPLIT 426 q850 q851
XSPLIT427 LSmitll_SPLIT 427 q852 q853
XSPLIT428 LSmitll_SPLIT 428 q854 q855
XSPLIT429 LSmitll_SPLIT 429 q856 q857
XSPLIT430 LSmitll_SPLIT 430 q858 q859
XSPLIT431 LSmitll_SPLIT 431 q860 q861
XSPLIT432 LSmitll_SPLIT 432 q862 q863
XSPLIT433 LSmitll_SPLIT 433 q864 q865
XSPLIT434 LSmitll_SPLIT 434 q866 q867
XSPLIT435 LSmitll_SPLIT 435 q868 q869
XSPLIT436 LSmitll_SPLIT 436 q870 q871
XSPLIT437 LSmitll_SPLIT 437 q872 q873
XSPLIT438 LSmitll_SPLIT 438 q874 q875
XSPLIT439 LSmitll_SPLIT 439 q876 q877
XSPLIT440 LSmitll_SPLIT 440 q878 q879
XSPLIT441 LSmitll_SPLIT 441 q880 q881
XSPLIT442 LSmitll_SPLIT 442 q882 q883
XSPLIT443 LSmitll_SPLIT 443 q884 q885
XSPLIT444 LSmitll_SPLIT 444 q886 q887
XSPLIT445 LSmitll_SPLIT 445 q888 q889
XSPLIT446 LSmitll_SPLIT 446 q890 q891
XSPLIT447 LSmitll_SPLIT 447 q892 q893
XSPLIT448 LSmitll_SPLIT 448 q894 q895
XSPLIT449 LSmitll_SPLIT 449 q896 q897
XSPLIT450 LSmitll_SPLIT 450 q898 q899
XSPLIT451 LSmitll_SPLIT 451 q900 q901
XSPLIT452 LSmitll_SPLIT 452 q902 q903
XSPLIT453 LSmitll_SPLIT 453 q904 q905
XSPLIT454 LSmitll_SPLIT 454 q906 q907
XSPLIT455 LSmitll_SPLIT 455 q908 q909
XSPLIT456 LSmitll_SPLIT 456 q910 q911
XSPLIT457 LSmitll_SPLIT 457 q912 q913
XSPLIT458 LSmitll_SPLIT 458 q914 q915
XSPLIT459 LSmitll_SPLIT 459 q916 q917
XSPLIT460 LSmitll_SPLIT 460 q918 q919
XSPLIT461 LSmitll_SPLIT 461 q920 q921
XSPLIT462 LSmitll_SPLIT 462 q922 q923
XSPLIT463 LSmitll_SPLIT 463 q924 q925
XSPLIT464 LSmitll_SPLIT 464 q926 q927
XSPLIT465 LSmitll_SPLIT 465 q928 q929
XSPLIT466 LSmitll_SPLIT 466 q930 q931
XSPLIT467 LSmitll_SPLIT 467 q932 q933
XSPLIT468 LSmitll_SPLIT 468 q934 q935
XSPLIT469 LSmitll_SPLIT 469 q936 q937
XSPLIT470 LSmitll_SPLIT 470 q938 q939
XSPLIT471 LSmitll_SPLIT 471 q940 q941
XSPLIT472 LSmitll_SPLIT 472 q942 q943
XSPLIT473 LSmitll_SPLIT 473 q944 q945
XSPLIT474 LSmitll_SPLIT 474 q946 q947
XSPLIT475 LSmitll_SPLIT 475 q948 q949
XSPLIT476 LSmitll_SPLIT 476 q950 q951
XSPLIT477 LSmitll_SPLIT 477 q952 q953
XSPLIT478 LSmitll_SPLIT 478 q954 q955
XSPLIT479 LSmitll_SPLIT 479 q956 q957
XSPLIT480 LSmitll_SPLIT 480 q958 q959
XSPLIT481 LSmitll_SPLIT 481 q960 q961
XSPLIT482 LSmitll_SPLIT 482 q962 q963
XSPLIT483 LSmitll_SPLIT 483 q964 q965
XSPLIT484 LSmitll_SPLIT 484 q966 q967
XSPLIT485 LSmitll_SPLIT 485 q968 q969
XSPLIT486 LSmitll_SPLIT 486 q970 q971
XSPLIT487 LSmitll_SPLIT 487 q972 q973
XSPLIT488 LSmitll_SPLIT 488 q974 q975
XSPLIT489 LSmitll_SPLIT 489 q976 q977
XSPLIT490 LSmitll_SPLIT 490 q978 q979
XSPLIT491 LSmitll_SPLIT 491 q980 q981
XSPLIT492 LSmitll_SPLIT 492 q982 q983
XSPLIT493 LSmitll_SPLIT 493 q984 q985
XSPLIT494 LSmitll_SPLIT 494 q986 q987
XSPLIT495 LSmitll_SPLIT 495 q988 q989
XSPLIT496 LSmitll_SPLIT 496 q990 q991
XSPLIT497 LSmitll_SPLIT 497 q992 q993
XSPLIT498 LSmitll_SPLIT 498 q994 q995
XSPLIT499 LSmitll_SPLIT 499 q996 q997
XSPLIT500 LSmitll_SPLIT 500 q998 q999
XSPLIT501 LSmitll_SPLIT 501 q1000 q1001
XSPLIT502 LSmitll_SPLIT 502 q1002 q1003
XSPLIT503 LSmitll_SPLIT 503 q1004 q1005
XSPLIT504 LSmitll_SPLIT 504 q1006 q1007
XSPLIT505 LSmitll_SPLIT 505 q1008 q1009
XSPLIT506 LSmitll_SPLIT 506 q1010 q1011
XSPLIT507 LSmitll_SPLIT 507 q1012 q1013
XSPLIT508 LSmitll_SPLIT 508 q1014 q1015
XSPLIT509 LSmitll_SPLIT 509 q1016 q1017
XSPLIT510 LSmitll_SPLIT 510 q1018 q1019
XSPLIT511 LSmitll_SPLIT 511 q1020 q1021
XSPLIT512 LSmitll_SPLIT 512 q1022 q1023
XSPLIT513 LSmitll_SPLIT 513 q1024 q1025
XSPLIT514 LSmitll_SPLIT 514 q1026 q1027
XSPLIT515 LSmitll_SPLIT 515 q1028 q1029
XSPLIT516 LSmitll_SPLIT 516 q1030 q1031
XSPLIT517 LSmitll_SPLIT 517 q1032 q1033
XSPLIT518 LSmitll_SPLIT 518 q1034 q1035
XSPLIT519 LSmitll_SPLIT 519 q1036 q1037
XSPLIT520 LSmitll_SPLIT 520 q1038 q1039
XSPLIT521 LSmitll_SPLIT 521 q1040 q1041
XSPLIT522 LSmitll_SPLIT 522 q1042 q1043
XSPLIT523 LSmitll_SPLIT 523 q1044 q1045
XSPLIT524 LSmitll_SPLIT 524 q1046 q1047
XSPLIT525 LSmitll_SPLIT 525 q1048 q1049
XSPLIT526 LSmitll_SPLIT 526 q1050 q1051
XSPLIT527 LSmitll_SPLIT 527 q1052 q1053
XSPLIT528 LSmitll_SPLIT 528 q1054 q1055
XSPLIT529 LSmitll_SPLIT 529 q1056 q1057
XSPLIT530 LSmitll_SPLIT 530 q1058 q1059
XSPLIT531 LSmitll_SPLIT 531 q1060 q1061
XSPLIT532 LSmitll_SPLIT 532 q1062 q1063
XSPLIT533 LSmitll_SPLIT 533 q1064 q1065
XSPLIT534 LSmitll_SPLIT 534 q1066 q1067
XSPLIT535 LSmitll_SPLIT 535 q1068 q1069
XSPLIT536 LSmitll_SPLIT 536 q1070 q1071
XSPLIT537 LSmitll_SPLIT 537 q1072 q1073
XSPLIT538 LSmitll_SPLIT 538 q1074 q1075
XSPLIT539 LSmitll_SPLIT 539 q1076 q1077
XSPLIT540 LSmitll_SPLIT 540 q1078 q1079
XSPLIT541 LSmitll_SPLIT 541 q1080 q1081
XSPLIT542 LSmitll_SPLIT 542 q1082 q1083
XSPLIT543 LSmitll_SPLIT 543 q1084 q1085
XSPLIT544 LSmitll_SPLIT 544 q1086 q1087
XSPLIT545 LSmitll_SPLIT 545 q1088 q1089
XSPLIT546 LSmitll_SPLIT 546 q1090 q1091
XSPLIT547 LSmitll_SPLIT 547 q1092 q1093
XSPLIT548 LSmitll_SPLIT 548 q1094 q1095
XSPLIT549 LSmitll_SPLIT 549 q1096 q1097
XSPLIT550 LSmitll_SPLIT 550 q1098 q1099
XSPLIT551 LSmitll_SPLIT 551 q1100 q1101
XSPLIT552 LSmitll_SPLIT 552 q1102 q1103
XSPLIT553 LSmitll_SPLIT 553 q1104 q1105
XSPLIT554 LSmitll_SPLIT 554 q1106 q1107
XSPLIT555 LSmitll_SPLIT 555 q1108 q1109
XSPLIT556 LSmitll_SPLIT 556 q1110 q1111
XSPLIT557 LSmitll_SPLIT 557 q1112 q1113
XSPLIT558 LSmitll_SPLIT 558 q1114 q1115
XSPLIT559 LSmitll_SPLIT 559 q1116 q1117
XSPLIT560 LSmitll_SPLIT 560 q1118 q1119
XSPLIT561 LSmitll_SPLIT 561 q1120 q1121
XSPLIT562 LSmitll_SPLIT 562 q1122 q1123
XSPLIT563 LSmitll_SPLIT 563 q1124 q1125
XSPLIT564 LSmitll_SPLIT 564 q1126 q1127
XSPLIT565 LSmitll_SPLIT 565 q1128 q1129
XSPLIT566 LSmitll_SPLIT 566 q1130 q1131
XSPLIT567 LSmitll_SPLIT 567 q1132 q1133
XSPLIT568 LSmitll_SPLIT 568 q1134 q1135
XSPLIT569 LSmitll_SPLIT 569 q1136 q1137
XSPLIT570 LSmitll_SPLIT 570 q1138 q1139
XSPLIT571 LSmitll_SPLIT 571 q1140 q1141
XSPLIT572 LSmitll_SPLIT 572 q1142 q1143
XSPLIT573 LSmitll_SPLIT 573 q1144 q1145
XSPLIT574 LSmitll_SPLIT 574 q1146 q1147
XSPLIT575 LSmitll_SPLIT 575 q1148 q1149
XSPLIT576 LSmitll_SPLIT 576 q1150 q1151
XSPLIT577 LSmitll_SPLIT 577 q1152 q1153
XSPLIT578 LSmitll_SPLIT 578 q1154 q1155
XSPLIT579 LSmitll_SPLIT 579 q1156 q1157
XSPLIT580 LSmitll_SPLIT 580 q1158 q1159
XSPLIT581 LSmitll_SPLIT 581 q1160 q1161
XSPLIT582 LSmitll_SPLIT 582 q1162 q1163
XSPLIT583 LSmitll_SPLIT 583 q1164 q1165
XSPLIT584 LSmitll_SPLIT 584 q1166 q1167
XSPLIT585 LSmitll_SPLIT 585 q1168 q1169
XSPLIT586 LSmitll_SPLIT 586 q1170 q1171
XSPLIT587 LSmitll_SPLIT 587 q1172 q1173
XSPLIT588 LSmitll_SPLIT 588 q1174 q1175
XSPLIT589 LSmitll_SPLIT 589 q1176 q1177
XSPLIT590 LSmitll_SPLIT 590 q1178 q1179
XSPLIT591 LSmitll_SPLIT 591 q1180 q1181
XSPLIT592 LSmitll_SPLIT 592 q1182 q1183
XSPLIT593 LSmitll_SPLIT 593 q1184 q1185
XSPLIT594 LSmitll_SPLIT 594 q1186 q1187
XSPLIT595 LSmitll_SPLIT 595 q1188 q1189
XSPLIT596 LSmitll_SPLIT 596 q1190 q1191
XSPLIT597 LSmitll_SPLIT 597 q1192 q1193
XSPLIT598 LSmitll_SPLIT 598 q1194 q1195
XSPLIT599 LSmitll_SPLIT 599 q1196 q1197
XSPLIT600 LSmitll_SPLIT 600 q1198 q1199
XSPLIT601 LSmitll_SPLIT 601 q1200 q1201
XSPLIT602 LSmitll_SPLIT 602 q1202 q1203
XSPLIT603 LSmitll_SPLIT 603 q1204 q1205
XSPLIT604 LSmitll_SPLIT 604 q1206 q1207
XSPLIT605 LSmitll_SPLIT 605 q1208 q1209
XSPLIT606 LSmitll_SPLIT 606 q1210 q1211
XSPLIT607 LSmitll_SPLIT 607 q1212 q1213
XSPLIT608 LSmitll_SPLIT 608 q1214 q1215
XSPLIT609 LSmitll_SPLIT 609 q1216 q1217
XSPLIT610 LSmitll_SPLIT 610 q1218 q1219
XSPLIT611 LSmitll_SPLIT 611 q1220 q1221
XSPLIT612 LSmitll_SPLIT 612 q1222 q1223
XSPLIT613 LSmitll_SPLIT 613 q1224 q1225
XSPLIT614 LSmitll_SPLIT 614 q1226 q1227
XSPLIT615 LSmitll_SPLIT 615 q1228 q1229
XSPLIT616 LSmitll_SPLIT 616 q1230 q1231
XSPLIT617 LSmitll_SPLIT 617 q1232 q1233
XSPLIT618 LSmitll_SPLIT 618 q1234 q1235
XSPLIT619 LSmitll_SPLIT 619 q1236 q1237
XSPLIT620 LSmitll_SPLIT 620 q1238 q1239
XSPLIT621 LSmitll_SPLIT 621 q1240 q1241
XSPLIT622 LSmitll_SPLIT 622 q1242 q1243
XSPLIT623 LSmitll_SPLIT 623 q1244 q1245
XSPLIT624 LSmitll_SPLIT 624 q1246 q1247
XSPLIT625 LSmitll_SPLIT 625 q1248 q1249
XSPLIT626 LSmitll_SPLIT 626 q1250 q1251
XSPLIT627 LSmitll_SPLIT 627 q1252 q1253
XSPLIT628 LSmitll_SPLIT 628 q1254 q1255
XSPLIT629 LSmitll_SPLIT 629 q1256 q1257
XSPLIT630 LSmitll_SPLIT 630 q1258 q1259
XSPLIT631 LSmitll_SPLIT 631 q1260 q1261
XSPLIT632 LSmitll_SPLIT 632 q1262 q1263
XSPLIT633 LSmitll_SPLIT 633 q1264 q1265
XSPLIT634 LSmitll_SPLIT 634 q1266 q1267
XSPLIT635 LSmitll_SPLIT 635 q1268 q1269
XSPLIT636 LSmitll_SPLIT 636 q1270 q1271
XSPLIT637 LSmitll_SPLIT 637 q1272 q1273
XSPLIT638 LSmitll_SPLIT 638 q1274 q1275
XSPLIT639 LSmitll_SPLIT 639 q1276 q1277
XSPLIT640 LSmitll_SPLIT 640 q1278 q1279
XSPLIT641 LSmitll_SPLIT 641 q1280 q1281
XSPLIT642 LSmitll_SPLIT 642 q1282 q1283
XSPLIT643 LSmitll_SPLIT 643 q1284 q1285
XSPLIT644 LSmitll_SPLIT 644 q1286 q1287
XSPLIT645 LSmitll_SPLIT 645 q1288 q1289
XSPLIT646 LSmitll_SPLIT 646 q1290 q1291
XSPLIT647 LSmitll_SPLIT 647 q1292 q1293
XSPLIT648 LSmitll_SPLIT 648 q1294 q1295
XSPLIT649 LSmitll_SPLIT 649 q1296 q1297
XSPLIT650 LSmitll_SPLIT 650 q1298 q1299
XSPLIT651 LSmitll_SPLIT 651 q1300 q1301
XSPLIT652 LSmitll_SPLIT 652 q1302 q1303
XSPLIT653 LSmitll_SPLIT 653 q1304 q1305
XSPLIT654 LSmitll_SPLIT 654 q1306 q1307
XSPLIT655 LSmitll_SPLIT 655 q1308 q1309
XSPLIT656 LSmitll_SPLIT 656 q1310 q1311
XSPLIT657 LSmitll_SPLIT 657 q1312 q1313
XSPLIT658 LSmitll_SPLIT 658 q1314 q1315
XSPLIT659 LSmitll_SPLIT 659 q1316 q1317
XSPLIT660 LSmitll_SPLIT 660 q1318 q1319
XSPLIT661 LSmitll_SPLIT 661 q1320 q1321
XSPLIT662 LSmitll_SPLIT 662 q1322 q1323
XSPLIT663 LSmitll_SPLIT 663 q1324 q1325
XSPLIT664 LSmitll_SPLIT 664 q1326 q1327
XSPLIT665 LSmitll_SPLIT 665 q1328 q1329
XSPLIT666 LSmitll_SPLIT 666 q1330 q1331
XSPLIT667 LSmitll_SPLIT 667 q1332 q1333
XSPLIT668 LSmitll_SPLIT 668 q1334 q1335
XSPLIT669 LSmitll_SPLIT 669 q1336 q1337
XSPLIT670 LSmitll_SPLIT 670 q1338 q1339
XSPLIT671 LSmitll_SPLIT 671 q1340 q1341
XSPLIT672 LSmitll_SPLIT 672 q1342 q1343
XSPLIT673 LSmitll_SPLIT 673 q1344 q1345
XSPLIT674 LSmitll_SPLIT 674 q1346 q1347
XSPLIT675 LSmitll_SPLIT 675 q1348 q1349
XSPLIT676 LSmitll_SPLIT 676 q1350 q1351
XSPLIT677 LSmitll_SPLIT 677 q1352 q1353
XSPLIT678 LSmitll_SPLIT 678 q1354 q1355
XSPLIT679 LSmitll_SPLIT 679 q1356 q1357
XSPLIT680 LSmitll_SPLIT 680 q1358 q1359
XSPLIT681 LSmitll_SPLIT 681 q1360 q1361
XSPLIT682 LSmitll_SPLIT 682 q1362 q1363
XSPLIT683 LSmitll_SPLIT 683 q1364 q1365
XSPLIT684 LSmitll_SPLIT 684 q1366 q1367
XSPLIT685 LSmitll_SPLIT 685 q1368 q1369
XSPLIT686 LSmitll_SPLIT 686 q1370 q1371
XSPLIT687 LSmitll_SPLIT 687 q1372 q1373
XSPLIT688 LSmitll_SPLIT 688 q1374 q1375
XSPLIT689 LSmitll_SPLIT 689 q1376 q1377
XSPLIT690 LSmitll_SPLIT 690 q1378 q1379
XSPLIT691 LSmitll_SPLIT 691 q1380 q1381
XSPLIT692 LSmitll_SPLIT 692 q1382 q1383
XSPLIT693 LSmitll_SPLIT 693 q1384 q1385
XSPLIT694 LSmitll_SPLIT 694 q1386 q1387
XSPLIT695 LSmitll_SPLIT 695 q1388 q1389
XSPLIT696 LSmitll_SPLIT 696 q1390 q1391
XSPLIT697 LSmitll_SPLIT 697 q1392 q1393
XSPLIT698 LSmitll_SPLIT 698 q1394 q1395
XSPLIT699 LSmitll_SPLIT 699 q1396 q1397
XSPLIT700 LSmitll_SPLIT 700 q1398 q1399
XSPLIT701 LSmitll_SPLIT 701 q1400 q1401
XSPLIT702 LSmitll_SPLIT 702 q1402 q1403
XSPLIT703 LSmitll_SPLIT 703 q1404 q1405
XSPLIT704 LSmitll_SPLIT 704 q1406 q1407
XSPLIT705 LSmitll_SPLIT 705 q1408 q1409
XSPLIT706 LSmitll_SPLIT 706 q1410 q1411
XSPLIT707 LSmitll_SPLIT 707 q1412 q1413
XSPLIT708 LSmitll_SPLIT 708 q1414 q1415
XSPLIT709 LSmitll_SPLIT 709 q1416 q1417
XSPLIT710 LSmitll_SPLIT 710 q1418 q1419
XSPLIT711 LSmitll_SPLIT 711 q1420 q1421
XSPLIT712 LSmitll_SPLIT 712 q1422 q1423
XSPLIT713 LSmitll_SPLIT 713 q1424 q1425
XSPLIT714 LSmitll_SPLIT 714 q1426 q1427
XSPLIT715 LSmitll_SPLIT 715 q1428 q1429
XSPLIT716 LSmitll_SPLIT 716 q1430 q1431
XSPLIT717 LSmitll_SPLIT 717 q1432 q1433
XSPLIT718 LSmitll_SPLIT 718 q1434 q1435
XSPLIT719 LSmitll_SPLIT 719 q1436 q1437
XSPLIT720 LSmitll_SPLIT 720 q1438 q1439
XSPLIT721 LSmitll_SPLIT 721 q1440 q1441
XSPLIT722 LSmitll_SPLIT 722 q1442 q1443
XSPLIT723 LSmitll_SPLIT 723 q1444 q1445
XSPLIT724 LSmitll_SPLIT 724 q1446 q1447
XSPLIT725 LSmitll_SPLIT 725 q1448 q1449
XSPLIT726 LSmitll_SPLIT 726 q1450 q1451
XSPLIT727 LSmitll_SPLIT 727 q1452 q1453
XSPLIT728 LSmitll_SPLIT 728 q1454 q1455
XSPLIT729 LSmitll_SPLIT 729 q1456 q1457
XSPLIT730 LSmitll_SPLIT 730 q1458 q1459
XSPLIT731 LSmitll_SPLIT 731 q1460 q1461
XSPLIT732 LSmitll_SPLIT 732 q1462 q1463
XSPLIT733 LSmitll_SPLIT 733 q1464 q1465
XSPLIT734 LSmitll_SPLIT 734 q1466 q1467
XSPLIT735 LSmitll_SPLIT 735 q1468 q1469
XSPLIT736 LSmitll_SPLIT 736 q1470 q1471
XSPLIT737 LSmitll_SPLIT 737 q1472 q1473
XSPLIT738 LSmitll_SPLIT 738 q1474 q1475
XSPLIT739 LSmitll_SPLIT 739 q1476 q1477
XSPLIT740 LSmitll_SPLIT 740 q1478 q1479
XSPLIT741 LSmitll_SPLIT 741 q1480 q1481
XSPLIT742 LSmitll_SPLIT 742 q1482 q1483
XSPLIT743 LSmitll_SPLIT 743 q1484 q1485
XSPLIT744 LSmitll_SPLIT 744 q1486 q1487
XSPLIT745 LSmitll_SPLIT 745 q1488 q1489
XSPLIT746 LSmitll_SPLIT 746 q1490 q1491
XSPLIT747 LSmitll_SPLIT 747 q1492 q1493
XSPLIT748 LSmitll_SPLIT 748 q1494 q1495
XSPLIT749 LSmitll_SPLIT 749 q1496 q1497
XSPLIT750 LSmitll_SPLIT 750 q1498 q1499
XSPLIT751 LSmitll_SPLIT 751 q1500 q1501
XSPLIT752 LSmitll_SPLIT 752 q1502 q1503
XSPLIT753 LSmitll_SPLIT 753 q1504 q1505
XSPLIT754 LSmitll_SPLIT 754 q1506 q1507
XSPLIT755 LSmitll_SPLIT 755 q1508 q1509
XSPLIT756 LSmitll_SPLIT 756 q1510 q1511
XSPLIT757 LSmitll_SPLIT 757 q1512 q1513
XSPLIT758 LSmitll_SPLIT 758 q1514 q1515
XSPLIT759 LSmitll_SPLIT 759 q1516 q1517
XSPLIT760 LSmitll_SPLIT 760 q1518 q1519
XSPLIT761 LSmitll_SPLIT 761 q1520 q1521
XSPLIT762 LSmitll_SPLIT 762 q1522 q1523
XSPLIT763 LSmitll_SPLIT 763 q1524 q1525
XSPLIT764 LSmitll_SPLIT 764 q1526 q1527
XSPLIT765 LSmitll_SPLIT 765 q1528 q1529
XSPLIT766 LSmitll_SPLIT 766 q1530 q1531
XSPLIT767 LSmitll_SPLIT 767 q1532 q1533
XSPLIT768 LSmitll_SPLIT 768 q1534 q1535
XSPLIT769 LSmitll_SPLIT 769 q1536 q1537
XSPLIT770 LSmitll_SPLIT 770 q1538 q1539
XSPLIT771 LSmitll_SPLIT 771 q1540 q1541
XSPLIT772 LSmitll_SPLIT 772 q1542 q1543
XSPLIT773 LSmitll_SPLIT 773 q1544 q1545
XSPLIT774 LSmitll_SPLIT 774 q1546 q1547
XSPLIT775 LSmitll_SPLIT 775 q1548 q1549
XSPLIT776 LSmitll_SPLIT 776 q1550 q1551
XSPLIT777 LSmitll_SPLIT 777 q1552 q1553
XSPLIT778 LSmitll_SPLIT 778 q1554 q1555
XSPLIT779 LSmitll_SPLIT 779 q1556 q1557
XSPLIT780 LSmitll_SPLIT 780 q1558 q1559
XSPLIT781 LSmitll_SPLIT 781 q1560 q1561
XSPLIT782 LSmitll_SPLIT 782 q1562 q1563
XSPLIT783 LSmitll_SPLIT 783 q1564 q1565
XSPLIT784 LSmitll_SPLIT 784 q1566 q1567
XSPLIT785 LSmitll_SPLIT 785 q1568 q1569
XSPLIT786 LSmitll_SPLIT 786 q1570 q1571
XSPLIT787 LSmitll_SPLIT 787 q1572 q1573
XSPLIT788 LSmitll_SPLIT 788 q1574 q1575
XSPLIT789 LSmitll_SPLIT 789 q1576 q1577
XSPLIT790 LSmitll_SPLIT 790 q1578 q1579
XSPLIT791 LSmitll_SPLIT 791 q1580 q1581
XSPLIT792 LSmitll_SPLIT 792 q1582 q1583
XSPLIT793 LSmitll_SPLIT 793 q1584 q1585
XSPLIT794 LSmitll_SPLIT 794 q1586 q1587
XSPLIT795 LSmitll_SPLIT 795 q1588 q1589
XSPLIT796 LSmitll_SPLIT 796 q1590 q1591
XSPLIT797 LSmitll_SPLIT 797 q1592 q1593
XSPLIT798 LSmitll_SPLIT 798 q1594 q1595
XSPLIT799 LSmitll_SPLIT 799 q1596 q1597
XSPLIT800 LSmitll_SPLIT 800 q1598 q1599
XSPLIT801 LSmitll_SPLIT 801 q1600 q1601
XSPLIT802 LSmitll_SPLIT 802 q1602 q1603
XSPLIT803 LSmitll_SPLIT 803 q1604 q1605
XSPLIT804 LSmitll_SPLIT 804 q1606 q1607
XSPLIT805 LSmitll_SPLIT 805 q1608 q1609
XSPLIT806 LSmitll_SPLIT 806 q1610 q1611
XSPLIT807 LSmitll_SPLIT 807 q1612 q1613
XSPLIT808 LSmitll_SPLIT 808 q1614 q1615
XSPLIT809 LSmitll_SPLIT 809 q1616 q1617
XSPLIT810 LSmitll_SPLIT 810 q1618 q1619
XSPLIT811 LSmitll_SPLIT 811 q1620 q1621
XSPLIT812 LSmitll_SPLIT 812 q1622 q1623
XSPLIT813 LSmitll_SPLIT 813 q1624 q1625
XSPLIT814 LSmitll_SPLIT 814 q1626 q1627
XSPLIT815 LSmitll_SPLIT 815 q1628 q1629
XSPLIT816 LSmitll_SPLIT 816 q1630 q1631
XSPLIT817 LSmitll_SPLIT 817 q1632 q1633
XSPLIT818 LSmitll_SPLIT 818 q1634 q1635
XSPLIT819 LSmitll_SPLIT 819 q1636 q1637
XSPLIT820 LSmitll_SPLIT 820 q1638 q1639
XSPLIT821 LSmitll_SPLIT 821 q1640 q1641
XSPLIT822 LSmitll_SPLIT 822 q1642 q1643
XSPLIT823 LSmitll_SPLIT 823 q1644 q1645
XSPLIT824 LSmitll_SPLIT 824 q1646 q1647
XSPLIT825 LSmitll_SPLIT 825 q1648 q1649
XSPLIT826 LSmitll_SPLIT 826 q1650 q1651
XSPLIT827 LSmitll_SPLIT 827 q1652 q1653
XSPLIT828 LSmitll_SPLIT 828 q1654 q1655
XSPLIT829 LSmitll_SPLIT 829 q1656 q1657
XSPLIT830 LSmitll_SPLIT 830 q1658 q1659
XSPLIT831 LSmitll_SPLIT 831 q1660 q1661
XSPLIT832 LSmitll_SPLIT 832 q1662 q1663
XSPLIT833 LSmitll_SPLIT 833 q1664 q1665
XSPLIT834 LSmitll_SPLIT 834 q1666 q1667
XSPLIT835 LSmitll_SPLIT 835 q1668 q1669
XSPLIT836 LSmitll_SPLIT 836 q1670 q1671
XSPLIT837 LSmitll_SPLIT 837 q1672 q1673
XSPLIT838 LSmitll_SPLIT 838 q1674 q1675
XSPLIT839 LSmitll_SPLIT 839 q1676 q1677
XSPLIT840 LSmitll_SPLIT 840 q1678 q1679
XSPLIT841 LSmitll_SPLIT 841 q1680 q1681
XSPLIT842 LSmitll_SPLIT 842 q1682 q1683
XSPLIT843 LSmitll_SPLIT 843 q1684 q1685
XSPLIT844 LSmitll_SPLIT 844 q1686 q1687
XSPLIT845 LSmitll_SPLIT 845 q1688 q1689
XSPLIT846 LSmitll_SPLIT 846 q1690 q1691
XSPLIT847 LSmitll_SPLIT 847 q1692 q1693
XSPLIT848 LSmitll_SPLIT 848 q1694 q1695
XSPLIT849 LSmitll_SPLIT 849 q1696 q1697
XSPLIT850 LSmitll_SPLIT 850 q1698 q1699
XSPLIT851 LSmitll_SPLIT 851 q1700 q1701
XSPLIT852 LSmitll_SPLIT 852 q1702 q1703
XSPLIT853 LSmitll_SPLIT 853 q1704 q1705
XSPLIT854 LSmitll_SPLIT 854 q1706 q1707
XSPLIT855 LSmitll_SPLIT 855 q1708 q1709
XSPLIT856 LSmitll_SPLIT 856 q1710 q1711
XSPLIT857 LSmitll_SPLIT 857 q1712 q1713
XSPLIT858 LSmitll_SPLIT 858 q1714 q1715
XSPLIT859 LSmitll_SPLIT 859 q1716 q1717
XSPLIT860 LSmitll_SPLIT 860 q1718 q1719
XSPLIT861 LSmitll_SPLIT 861 q1720 q1721
XSPLIT862 LSmitll_SPLIT 862 q1722 q1723
XSPLIT863 LSmitll_SPLIT 863 q1724 q1725
XSPLIT864 LSmitll_SPLIT 864 q1726 q1727
XSPLIT865 LSmitll_SPLIT 865 q1728 q1729
XSPLIT866 LSmitll_SPLIT 866 q1730 q1731
XSPLIT867 LSmitll_SPLIT 867 q1732 q1733
XSPLIT868 LSmitll_SPLIT 868 q1734 q1735
XSPLIT869 LSmitll_SPLIT 869 q1736 q1737
XSPLIT870 LSmitll_SPLIT 870 q1738 q1739
XSPLIT871 LSmitll_SPLIT 871 q1740 q1741
XSPLIT872 LSmitll_SPLIT 872 q1742 q1743
XSPLIT873 LSmitll_SPLIT 873 q1744 q1745
XSPLIT874 LSmitll_SPLIT 874 q1746 q1747
XSPLIT875 LSmitll_SPLIT 875 q1748 q1749
XSPLIT876 LSmitll_SPLIT 876 q1750 q1751
XSPLIT877 LSmitll_SPLIT 877 q1752 q1753
XSPLIT878 LSmitll_SPLIT 878 q1754 q1755
XSPLIT879 LSmitll_SPLIT 879 q1756 q1757
XSPLIT880 LSmitll_SPLIT 880 q1758 q1759
XSPLIT881 LSmitll_SPLIT 881 q1760 q1761
XSPLIT882 LSmitll_SPLIT 882 q1762 q1763
XSPLIT883 LSmitll_SPLIT 883 q1764 q1765
XSPLIT884 LSmitll_SPLIT 884 q1766 q1767
XSPLIT885 LSmitll_SPLIT 885 q1768 q1769
XSPLIT886 LSmitll_SPLIT 886 q1770 q1771
XSPLIT887 LSmitll_SPLIT 887 q1772 q1773
XSPLIT888 LSmitll_SPLIT 888 q1774 q1775
XSPLIT889 LSmitll_SPLIT 889 q1776 q1777
XSPLIT890 LSmitll_SPLIT 890 q1778 q1779
XSPLIT891 LSmitll_SPLIT 891 q1780 q1781
XSPLIT892 LSmitll_SPLIT 892 q1782 q1783
XSPLIT893 LSmitll_SPLIT 893 q1784 q1785
XSPLIT894 LSmitll_SPLIT 894 q1786 q1787
XSPLIT895 LSmitll_SPLIT 895 q1788 q1789
XSPLIT896 LSmitll_SPLIT 896 q1790 q1791
XSPLIT897 LSmitll_SPLIT 897 q1792 q1793
XSPLIT898 LSmitll_SPLIT 898 q1794 q1795
XSPLIT899 LSmitll_SPLIT 899 q1796 q1797
XSPLIT900 LSmitll_SPLIT 900 q1798 q1799
XSPLIT901 LSmitll_SPLIT 901 q1800 q1801
XSPLIT902 LSmitll_SPLIT 902 q1802 q1803
XSPLIT903 LSmitll_SPLIT 903 q1804 q1805
XSPLIT904 LSmitll_SPLIT 904 q1806 q1807
XSPLIT905 LSmitll_SPLIT 905 q1808 q1809
XSPLIT906 LSmitll_SPLIT 906 q1810 q1811
XSPLIT907 LSmitll_SPLIT 907 q1812 q1813
XSPLIT908 LSmitll_SPLIT 908 q1814 q1815
XSPLIT909 LSmitll_SPLIT 909 q1816 q1817
XSPLIT910 LSmitll_SPLIT 910 q1818 q1819
XSPLIT911 LSmitll_SPLIT 911 q1820 q1821
XSPLIT912 LSmitll_SPLIT 912 q1822 q1823
XSPLIT913 LSmitll_SPLIT 913 q1824 q1825
XSPLIT914 LSmitll_SPLIT 914 q1826 q1827
XSPLIT915 LSmitll_SPLIT 915 q1828 q1829
XSPLIT916 LSmitll_SPLIT 916 q1830 q1831
XSPLIT917 LSmitll_SPLIT 917 q1832 q1833
XSPLIT918 LSmitll_SPLIT 918 q1834 q1835
XSPLIT919 LSmitll_SPLIT 919 q1836 q1837
XSPLIT920 LSmitll_SPLIT 920 q1838 q1839
XSPLIT921 LSmitll_SPLIT 921 q1840 q1841
XSPLIT922 LSmitll_SPLIT 922 q1842 q1843
XSPLIT923 LSmitll_SPLIT 923 q1844 q1845
XSPLIT924 LSmitll_SPLIT 924 q1846 q1847
XSPLIT925 LSmitll_SPLIT 925 q1848 q1849
XSPLIT926 LSmitll_SPLIT 926 q1850 q1851
XSPLIT927 LSmitll_SPLIT 927 q1852 q1853
XSPLIT928 LSmitll_SPLIT 928 q1854 q1855
XSPLIT929 LSmitll_SPLIT 929 q1856 q1857
XSPLIT930 LSmitll_SPLIT 930 q1858 q1859
XSPLIT931 LSmitll_SPLIT 931 q1860 q1861
XSPLIT932 LSmitll_SPLIT 932 q1862 q1863
XSPLIT933 LSmitll_SPLIT 933 q1864 q1865
XSPLIT934 LSmitll_SPLIT 934 q1866 q1867
XSPLIT935 LSmitll_SPLIT 935 q1868 q1869
XSPLIT936 LSmitll_SPLIT 936 q1870 q1871
XSPLIT937 LSmitll_SPLIT 937 q1872 q1873
XSPLIT938 LSmitll_SPLIT 938 q1874 q1875
XSPLIT939 LSmitll_SPLIT 939 q1876 q1877
XSPLIT940 LSmitll_SPLIT 940 q1878 q1879
XSPLIT941 LSmitll_SPLIT 941 q1880 q1881
XSPLIT942 LSmitll_SPLIT 942 q1882 q1883
XSPLIT943 LSmitll_SPLIT 943 q1884 q1885
XSPLIT944 LSmitll_SPLIT 944 q1886 q1887
XSPLIT945 LSmitll_SPLIT 945 q1888 q1889
XSPLIT946 LSmitll_SPLIT 946 q1890 q1891
XSPLIT947 LSmitll_SPLIT 947 q1892 q1893
XSPLIT948 LSmitll_SPLIT 948 q1894 q1895
XSPLIT949 LSmitll_SPLIT 949 q1896 q1897
XSPLIT950 LSmitll_SPLIT 950 q1898 q1899
XSPLIT951 LSmitll_SPLIT 951 q1900 q1901
XSPLIT952 LSmitll_SPLIT 952 q1902 q1903
XSPLIT953 LSmitll_SPLIT 953 q1904 q1905
XSPLIT954 LSmitll_SPLIT 954 q1906 q1907
XSPLIT955 LSmitll_SPLIT 955 q1908 q1909
XSPLIT956 LSmitll_SPLIT 956 q1910 q1911
XSPLIT957 LSmitll_SPLIT 957 q1912 q1913
XSPLIT958 LSmitll_SPLIT 958 q1914 q1915
XSPLIT959 LSmitll_SPLIT 959 q1916 q1917
XSPLIT960 LSmitll_SPLIT 960 q1918 q1919
XSPLIT961 LSmitll_SPLIT 961 q1920 q1921
XSPLIT962 LSmitll_SPLIT 962 q1922 q1923
XSPLIT963 LSmitll_SPLIT 963 q1924 q1925
XSPLIT964 LSmitll_SPLIT 964 q1926 q1927
XSPLIT965 LSmitll_SPLIT 965 q1928 q1929
XSPLIT966 LSmitll_SPLIT 966 q1930 q1931
XSPLIT967 LSmitll_SPLIT 967 q1932 q1933
XSPLIT968 LSmitll_SPLIT 968 q1934 q1935
XSPLIT969 LSmitll_SPLIT 969 q1936 q1937
XSPLIT970 LSmitll_SPLIT 970 q1938 q1939
XSPLIT971 LSmitll_SPLIT 971 q1940 q1941
XSPLIT972 LSmitll_SPLIT 972 q1942 q1943
XSPLIT973 LSmitll_SPLIT 973 q1944 q1945
XSPLIT974 LSmitll_SPLIT 974 q1946 q1947
XSPLIT975 LSmitll_SPLIT 975 q1948 q1949
XSPLIT976 LSmitll_SPLIT 976 q1950 q1951
XSPLIT977 LSmitll_SPLIT 977 q1952 q1953
XSPLIT978 LSmitll_SPLIT 978 q1954 q1955
XSPLIT979 LSmitll_SPLIT 979 q1956 q1957
XSPLIT980 LSmitll_SPLIT 980 q1958 q1959
XSPLIT981 LSmitll_SPLIT 981 q1960 q1961
XSPLIT982 LSmitll_SPLIT 982 q1962 q1963
XSPLIT983 LSmitll_SPLIT 983 q1964 q1965
XSPLIT984 LSmitll_SPLIT 984 q1966 q1967
XSPLIT985 LSmitll_SPLIT 985 q1968 q1969
XSPLIT986 LSmitll_SPLIT 986 q1970 q1971
XSPLIT987 LSmitll_SPLIT 987 q1972 q1973
XSPLIT988 LSmitll_SPLIT 988 q1974 q1975
XSPLIT989 LSmitll_SPLIT 989 q1976 q1977
XSPLIT990 LSmitll_SPLIT 990 q1978 q1979
XSPLIT991 LSmitll_SPLIT 991 q1980 q1981
XSPLIT992 LSmitll_SPLIT 992 q1982 q1983
XSPLIT993 LSmitll_SPLIT 993 q1984 q1985
XSPLIT994 LSmitll_SPLIT 994 q1986 q1987
XSPLIT995 LSmitll_SPLIT 995 q1988 q1989
XSPLIT996 LSmitll_SPLIT 996 q1990 q1991
XSPLIT997 LSmitll_SPLIT 997 q1992 q1993
XSPLIT998 LSmitll_SPLIT 998 q1994 q1995
XSPLIT999 LSmitll_SPLIT 999 q1996 q1997
XSPLIT1000 LSmitll_SPLIT 1000 q1998 q1999
XSPLIT1001 LSmitll_SPLIT 1001 q2000 q2001
XSPLIT1002 LSmitll_SPLIT 1002 q2002 q2003
XSPLIT1003 LSmitll_SPLIT 1003 q2004 q2005
XSPLIT1004 LSmitll_SPLIT 1004 q2006 q2007
XSPLIT1005 LSmitll_SPLIT 1005 q2008 q2009
XSPLIT1006 LSmitll_SPLIT 1006 q2010 q2011
XSPLIT1007 LSmitll_SPLIT 1007 q2012 q2013
XSPLIT1008 LSmitll_SPLIT 1008 q2014 q2015
XSPLIT1009 LSmitll_SPLIT 1009 q2016 q2017
XSPLIT1010 LSmitll_SPLIT 1010 q2018 q2019
XSPLIT1011 LSmitll_SPLIT 1011 q2020 q2021
XSPLIT1012 LSmitll_SPLIT 1012 q2022 q2023
XSPLIT1013 LSmitll_SPLIT 1013 q2024 q2025
XSPLIT1014 LSmitll_SPLIT 1014 q2026 q2027
XSPLIT1015 LSmitll_SPLIT 1015 q2028 q2029
XSPLIT1016 LSmitll_SPLIT 1016 q2030 q2031
XSPLIT1017 LSmitll_SPLIT 1017 q2032 q2033
XSPLIT1018 LSmitll_SPLIT 1018 q2034 q2035
XSPLIT1019 LSmitll_SPLIT 1019 q2036 q2037
XSPLIT1020 LSmitll_SPLIT 1020 q2038 q2039
XSPLIT1021 LSmitll_SPLIT 1021 q2040 q2041
XSPLIT1022 LSmitll_SPLIT 1022 q2042 q2043
XSPLIT1023 LSmitll_SPLIT 1023 q2044 q2045
XSPLIT1024 LSmitll_SPLIT 1024 q2046 q2047
.ends 1_to_2048_split

.subckt 1_to_1695_split a q0 q1 q2 q3 q4 q5 q6 q7 q8 q9 q10 q11 q12 q13 q14 q15 q16 q17 q18 q19 q20 q21 q22 q23 q24 q25 q26 q27 q28 q29 q30 q31 q32 q33 q34 q35 q36 q37 q38 q39 q40 q41 q42 q43 q44 q45 q46 q47 q48 q49 q50 q51 q52 q53 q54 q55 q56 q57 q58 q59 q60 q61 q62 q63 q64 q65 q66 q67 q68 q69 q70 q71 q72 q73 q74 q75 q76 q77 q78 q79 q80 q81 q82 q83 q84 q85 q86 q87 q88 q89 q90 q91 q92 q93 q94 q95 q96 q97 q98 q99 q100 q101 q102 q103 q104 q105 q106 q107 q108 q109 q110 q111 q112 q113 q114 q115 q116 q117 q118 q119 q120 q121 q122 q123 q124 q125 q126 q127 q128 q129 q130 q131 q132 q133 q134 q135 q136 q137 q138 q139 q140 q141 q142 q143 q144 q145 q146 q147 q148 q149 q150 q151 q152 q153 q154 q155 q156 q157 q158 q159 q160 q161 q162 q163 q164 q165 q166 q167 q168 q169 q170 q171 q172 q173 q174 q175 q176 q177 q178 q179 q180 q181 q182 q183 q184 q185 q186 q187 q188 q189 q190 q191 q192 q193 q194 q195 q196 q197 q198 q199 q200 q201 q202 q203 q204 q205 q206 q207 q208 q209 q210 q211 q212 q213 q214 q215 q216 q217 q218 q219 q220 q221 q222 q223 q224 q225 q226 q227 q228 q229 q230 q231 q232 q233 q234 q235 q236 q237 q238 q239 q240 q241 q242 q243 q244 q245 q246 q247 q248 q249 q250 q251 q252 q253 q254 q255 q256 q257 q258 q259 q260 q261 q262 q263 q264 q265 q266 q267 q268 q269 q270 q271 q272 q273 q274 q275 q276 q277 q278 q279 q280 q281 q282 q283 q284 q285 q286 q287 q288 q289 q290 q291 q292 q293 q294 q295 q296 q297 q298 q299 q300 q301 q302 q303 q304 q305 q306 q307 q308 q309 q310 q311 q312 q313 q314 q315 q316 q317 q318 q319 q320 q321 q322 q323 q324 q325 q326 q327 q328 q329 q330 q331 q332 q333 q334 q335 q336 q337 q338 q339 q340 q341 q342 q343 q344 q345 q346 q347 q348 q349 q350 q351 q352 q353 q354 q355 q356 q357 q358 q359 q360 q361 q362 q363 q364 q365 q366 q367 q368 q369 q370 q371 q372 q373 q374 q375 q376 q377 q378 q379 q380 q381 q382 q383 q384 q385 q386 q387 q388 q389 q390 q391 q392 q393 q394 q395 q396 q397 q398 q399 q400 q401 q402 q403 q404 q405 q406 q407 q408 q409 q410 q411 q412 q413 q414 q415 q416 q417 q418 q419 q420 q421 q422 q423 q424 q425 q426 q427 q428 q429 q430 q431 q432 q433 q434 q435 q436 q437 q438 q439 q440 q441 q442 q443 q444 q445 q446 q447 q448 q449 q450 q451 q452 q453 q454 q455 q456 q457 q458 q459 q460 q461 q462 q463 q464 q465 q466 q467 q468 q469 q470 q471 q472 q473 q474 q475 q476 q477 q478 q479 q480 q481 q482 q483 q484 q485 q486 q487 q488 q489 q490 q491 q492 q493 q494 q495 q496 q497 q498 q499 q500 q501 q502 q503 q504 q505 q506 q507 q508 q509 q510 q511 q512 q513 q514 q515 q516 q517 q518 q519 q520 q521 q522 q523 q524 q525 q526 q527 q528 q529 q530 q531 q532 q533 q534 q535 q536 q537 q538 q539 q540 q541 q542 q543 q544 q545 q546 q547 q548 q549 q550 q551 q552 q553 q554 q555 q556 q557 q558 q559 q560 q561 q562 q563 q564 q565 q566 q567 q568 q569 q570 q571 q572 q573 q574 q575 q576 q577 q578 q579 q580 q581 q582 q583 q584 q585 q586 q587 q588 q589 q590 q591 q592 q593 q594 q595 q596 q597 q598 q599 q600 q601 q602 q603 q604 q605 q606 q607 q608 q609 q610 q611 q612 q613 q614 q615 q616 q617 q618 q619 q620 q621 q622 q623 q624 q625 q626 q627 q628 q629 q630 q631 q632 q633 q634 q635 q636 q637 q638 q639 q640 q641 q642 q643 q644 q645 q646 q647 q648 q649 q650 q651 q652 q653 q654 q655 q656 q657 q658 q659 q660 q661 q662 q663 q664 q665 q666 q667 q668 q669 q670 q671 q672 q673 q674 q675 q676 q677 q678 q679 q680 q681 q682 q683 q684 q685 q686 q687 q688 q689 q690 q691 q692 q693 q694 q695 q696 q697 q698 q699 q700 q701 q702 q703 q704 q705 q706 q707 q708 q709 q710 q711 q712 q713 q714 q715 q716 q717 q718 q719 q720 q721 q722 q723 q724 q725 q726 q727 q728 q729 q730 q731 q732 q733 q734 q735 q736 q737 q738 q739 q740 q741 q742 q743 q744 q745 q746 q747 q748 q749 q750 q751 q752 q753 q754 q755 q756 q757 q758 q759 q760 q761 q762 q763 q764 q765 q766 q767 q768 q769 q770 q771 q772 q773 q774 q775 q776 q777 q778 q779 q780 q781 q782 q783 q784 q785 q786 q787 q788 q789 q790 q791 q792 q793 q794 q795 q796 q797 q798 q799 q800 q801 q802 q803 q804 q805 q806 q807 q808 q809 q810 q811 q812 q813 q814 q815 q816 q817 q818 q819 q820 q821 q822 q823 q824 q825 q826 q827 q828 q829 q830 q831 q832 q833 q834 q835 q836 q837 q838 q839 q840 q841 q842 q843 q844 q845 q846 q847 q848 q849 q850 q851 q852 q853 q854 q855 q856 q857 q858 q859 q860 q861 q862 q863 q864 q865 q866 q867 q868 q869 q870 q871 q872 q873 q874 q875 q876 q877 q878 q879 q880 q881 q882 q883 q884 q885 q886 q887 q888 q889 q890 q891 q892 q893 q894 q895 q896 q897 q898 q899 q900 q901 q902 q903 q904 q905 q906 q907 q908 q909 q910 q911 q912 q913 q914 q915 q916 q917 q918 q919 q920 q921 q922 q923 q924 q925 q926 q927 q928 q929 q930 q931 q932 q933 q934 q935 q936 q937 q938 q939 q940 q941 q942 q943 q944 q945 q946 q947 q948 q949 q950 q951 q952 q953 q954 q955 q956 q957 q958 q959 q960 q961 q962 q963 q964 q965 q966 q967 q968 q969 q970 q971 q972 q973 q974 q975 q976 q977 q978 q979 q980 q981 q982 q983 q984 q985 q986 q987 q988 q989 q990 q991 q992 q993 q994 q995 q996 q997 q998 q999 q1000 q1001 q1002 q1003 q1004 q1005 q1006 q1007 q1008 q1009 q1010 q1011 q1012 q1013 q1014 q1015 q1016 q1017 q1018 q1019 q1020 q1021 q1022 q1023 q1024 q1025 q1026 q1027 q1028 q1029 q1030 q1031 q1032 q1033 q1034 q1035 q1036 q1037 q1038 q1039 q1040 q1041 q1042 q1043 q1044 q1045 q1046 q1047 q1048 q1049 q1050 q1051 q1052 q1053 q1054 q1055 q1056 q1057 q1058 q1059 q1060 q1061 q1062 q1063 q1064 q1065 q1066 q1067 q1068 q1069 q1070 q1071 q1072 q1073 q1074 q1075 q1076 q1077 q1078 q1079 q1080 q1081 q1082 q1083 q1084 q1085 q1086 q1087 q1088 q1089 q1090 q1091 q1092 q1093 q1094 q1095 q1096 q1097 q1098 q1099 q1100 q1101 q1102 q1103 q1104 q1105 q1106 q1107 q1108 q1109 q1110 q1111 q1112 q1113 q1114 q1115 q1116 q1117 q1118 q1119 q1120 q1121 q1122 q1123 q1124 q1125 q1126 q1127 q1128 q1129 q1130 q1131 q1132 q1133 q1134 q1135 q1136 q1137 q1138 q1139 q1140 q1141 q1142 q1143 q1144 q1145 q1146 q1147 q1148 q1149 q1150 q1151 q1152 q1153 q1154 q1155 q1156 q1157 q1158 q1159 q1160 q1161 q1162 q1163 q1164 q1165 q1166 q1167 q1168 q1169 q1170 q1171 q1172 q1173 q1174 q1175 q1176 q1177 q1178 q1179 q1180 q1181 q1182 q1183 q1184 q1185 q1186 q1187 q1188 q1189 q1190 q1191 q1192 q1193 q1194 q1195 q1196 q1197 q1198 q1199 q1200 q1201 q1202 q1203 q1204 q1205 q1206 q1207 q1208 q1209 q1210 q1211 q1212 q1213 q1214 q1215 q1216 q1217 q1218 q1219 q1220 q1221 q1222 q1223 q1224 q1225 q1226 q1227 q1228 q1229 q1230 q1231 q1232 q1233 q1234 q1235 q1236 q1237 q1238 q1239 q1240 q1241 q1242 q1243 q1244 q1245 q1246 q1247 q1248 q1249 q1250 q1251 q1252 q1253 q1254 q1255 q1256 q1257 q1258 q1259 q1260 q1261 q1262 q1263 q1264 q1265 q1266 q1267 q1268 q1269 q1270 q1271 q1272 q1273 q1274 q1275 q1276 q1277 q1278 q1279 q1280 q1281 q1282 q1283 q1284 q1285 q1286 q1287 q1288 q1289 q1290 q1291 q1292 q1293 q1294 q1295 q1296 q1297 q1298 q1299 q1300 q1301 q1302 q1303 q1304 q1305 q1306 q1307 q1308 q1309 q1310 q1311 q1312 q1313 q1314 q1315 q1316 q1317 q1318 q1319 q1320 q1321 q1322 q1323 q1324 q1325 q1326 q1327 q1328 q1329 q1330 q1331 q1332 q1333 q1334 q1335 q1336 q1337 q1338 q1339 q1340 q1341 q1342 q1343 q1344 q1345 q1346 q1347 q1348 q1349 q1350 q1351 q1352 q1353 q1354 q1355 q1356 q1357 q1358 q1359 q1360 q1361 q1362 q1363 q1364 q1365 q1366 q1367 q1368 q1369 q1370 q1371 q1372 q1373 q1374 q1375 q1376 q1377 q1378 q1379 q1380 q1381 q1382 q1383 q1384 q1385 q1386 q1387 q1388 q1389 q1390 q1391 q1392 q1393 q1394 q1395 q1396 q1397 q1398 q1399 q1400 q1401 q1402 q1403 q1404 q1405 q1406 q1407 q1408 q1409 q1410 q1411 q1412 q1413 q1414 q1415 q1416 q1417 q1418 q1419 q1420 q1421 q1422 q1423 q1424 q1425 q1426 q1427 q1428 q1429 q1430 q1431 q1432 q1433 q1434 q1435 q1436 q1437 q1438 q1439 q1440 q1441 q1442 q1443 q1444 q1445 q1446 q1447 q1448 q1449 q1450 q1451 q1452 q1453 q1454 q1455 q1456 q1457 q1458 q1459 q1460 q1461 q1462 q1463 q1464 q1465 q1466 q1467 q1468 q1469 q1470 q1471 q1472 q1473 q1474 q1475 q1476 q1477 q1478 q1479 q1480 q1481 q1482 q1483 q1484 q1485 q1486 q1487 q1488 q1489 q1490 q1491 q1492 q1493 q1494 q1495 q1496 q1497 q1498 q1499 q1500 q1501 q1502 q1503 q1504 q1505 q1506 q1507 q1508 q1509 q1510 q1511 q1512 q1513 q1514 q1515 q1516 q1517 q1518 q1519 q1520 q1521 q1522 q1523 q1524 q1525 q1526 q1527 q1528 q1529 q1530 q1531 q1532 q1533 q1534 q1535 q1536 q1537 q1538 q1539 q1540 q1541 q1542 q1543 q1544 q1545 q1546 q1547 q1548 q1549 q1550 q1551 q1552 q1553 q1554 q1555 q1556 q1557 q1558 q1559 q1560 q1561 q1562 q1563 q1564 q1565 q1566 q1567 q1568 q1569 q1570 q1571 q1572 q1573 q1574 q1575 q1576 q1577 q1578 q1579 q1580 q1581 q1582 q1583 q1584 q1585 q1586 q1587 q1588 q1589 q1590 q1591 q1592 q1593 q1594 q1595 q1596 q1597 q1598 q1599 q1600 q1601 q1602 q1603 q1604 q1605 q1606 q1607 q1608 q1609 q1610 q1611 q1612 q1613 q1614 q1615 q1616 q1617 q1618 q1619 q1620 q1621 q1622 q1623 q1624 q1625 q1626 q1627 q1628 q1629 q1630 q1631 q1632 q1633 q1634 q1635 q1636 q1637 q1638 q1639 q1640 q1641 q1642 q1643 q1644 q1645 q1646 q1647 q1648 q1649 q1650 q1651 q1652 q1653 q1654 q1655 q1656 q1657 q1658 q1659 q1660 q1661 q1662 q1663 q1664 q1665 q1666 q1667 q1668 q1669 q1670 q1671 q1672 q1673 q1674 q1675 q1676 q1677 q1678 q1679 q1680 q1681 q1682 q1683 q1684 q1685 q1686 q1687 q1688 q1689 q1690 q1691 q1692 q1693 q1694 q1695 
XSPLIT_848 1_to_848_split a 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848
XSPLIT1 LSmitll_SPLIT 1 q0 q1
XSPLIT2 LSmitll_SPLIT 2 q2 q3
XSPLIT3 LSmitll_SPLIT 3 q4 q5
XSPLIT4 LSmitll_SPLIT 4 q6 q7
XSPLIT5 LSmitll_SPLIT 5 q8 q9
XSPLIT6 LSmitll_SPLIT 6 q10 q11
XSPLIT7 LSmitll_SPLIT 7 q12 q13
XSPLIT8 LSmitll_SPLIT 8 q14 q15
XSPLIT9 LSmitll_SPLIT 9 q16 q17
XSPLIT10 LSmitll_SPLIT 10 q18 q19
XSPLIT11 LSmitll_SPLIT 11 q20 q21
XSPLIT12 LSmitll_SPLIT 12 q22 q23
XSPLIT13 LSmitll_SPLIT 13 q24 q25
XSPLIT14 LSmitll_SPLIT 14 q26 q27
XSPLIT15 LSmitll_SPLIT 15 q28 q29
XSPLIT16 LSmitll_SPLIT 16 q30 q31
XSPLIT17 LSmitll_SPLIT 17 q32 q33
XSPLIT18 LSmitll_SPLIT 18 q34 q35
XSPLIT19 LSmitll_SPLIT 19 q36 q37
XSPLIT20 LSmitll_SPLIT 20 q38 q39
XSPLIT21 LSmitll_SPLIT 21 q40 q41
XSPLIT22 LSmitll_SPLIT 22 q42 q43
XSPLIT23 LSmitll_SPLIT 23 q44 q45
XSPLIT24 LSmitll_SPLIT 24 q46 q47
XSPLIT25 LSmitll_SPLIT 25 q48 q49
XSPLIT26 LSmitll_SPLIT 26 q50 q51
XSPLIT27 LSmitll_SPLIT 27 q52 q53
XSPLIT28 LSmitll_SPLIT 28 q54 q55
XSPLIT29 LSmitll_SPLIT 29 q56 q57
XSPLIT30 LSmitll_SPLIT 30 q58 q59
XSPLIT31 LSmitll_SPLIT 31 q60 q61
XSPLIT32 LSmitll_SPLIT 32 q62 q63
XSPLIT33 LSmitll_SPLIT 33 q64 q65
XSPLIT34 LSmitll_SPLIT 34 q66 q67
XSPLIT35 LSmitll_SPLIT 35 q68 q69
XSPLIT36 LSmitll_SPLIT 36 q70 q71
XSPLIT37 LSmitll_SPLIT 37 q72 q73
XSPLIT38 LSmitll_SPLIT 38 q74 q75
XSPLIT39 LSmitll_SPLIT 39 q76 q77
XSPLIT40 LSmitll_SPLIT 40 q78 q79
XSPLIT41 LSmitll_SPLIT 41 q80 q81
XSPLIT42 LSmitll_SPLIT 42 q82 q83
XSPLIT43 LSmitll_SPLIT 43 q84 q85
XSPLIT44 LSmitll_SPLIT 44 q86 q87
XSPLIT45 LSmitll_SPLIT 45 q88 q89
XSPLIT46 LSmitll_SPLIT 46 q90 q91
XSPLIT47 LSmitll_SPLIT 47 q92 q93
XSPLIT48 LSmitll_SPLIT 48 q94 q95
XSPLIT49 LSmitll_SPLIT 49 q96 q97
XSPLIT50 LSmitll_SPLIT 50 q98 q99
XSPLIT51 LSmitll_SPLIT 51 q100 q101
XSPLIT52 LSmitll_SPLIT 52 q102 q103
XSPLIT53 LSmitll_SPLIT 53 q104 q105
XSPLIT54 LSmitll_SPLIT 54 q106 q107
XSPLIT55 LSmitll_SPLIT 55 q108 q109
XSPLIT56 LSmitll_SPLIT 56 q110 q111
XSPLIT57 LSmitll_SPLIT 57 q112 q113
XSPLIT58 LSmitll_SPLIT 58 q114 q115
XSPLIT59 LSmitll_SPLIT 59 q116 q117
XSPLIT60 LSmitll_SPLIT 60 q118 q119
XSPLIT61 LSmitll_SPLIT 61 q120 q121
XSPLIT62 LSmitll_SPLIT 62 q122 q123
XSPLIT63 LSmitll_SPLIT 63 q124 q125
XSPLIT64 LSmitll_SPLIT 64 q126 q127
XSPLIT65 LSmitll_SPLIT 65 q128 q129
XSPLIT66 LSmitll_SPLIT 66 q130 q131
XSPLIT67 LSmitll_SPLIT 67 q132 q133
XSPLIT68 LSmitll_SPLIT 68 q134 q135
XSPLIT69 LSmitll_SPLIT 69 q136 q137
XSPLIT70 LSmitll_SPLIT 70 q138 q139
XSPLIT71 LSmitll_SPLIT 71 q140 q141
XSPLIT72 LSmitll_SPLIT 72 q142 q143
XSPLIT73 LSmitll_SPLIT 73 q144 q145
XSPLIT74 LSmitll_SPLIT 74 q146 q147
XSPLIT75 LSmitll_SPLIT 75 q148 q149
XSPLIT76 LSmitll_SPLIT 76 q150 q151
XSPLIT77 LSmitll_SPLIT 77 q152 q153
XSPLIT78 LSmitll_SPLIT 78 q154 q155
XSPLIT79 LSmitll_SPLIT 79 q156 q157
XSPLIT80 LSmitll_SPLIT 80 q158 q159
XSPLIT81 LSmitll_SPLIT 81 q160 q161
XSPLIT82 LSmitll_SPLIT 82 q162 q163
XSPLIT83 LSmitll_SPLIT 83 q164 q165
XSPLIT84 LSmitll_SPLIT 84 q166 q167
XSPLIT85 LSmitll_SPLIT 85 q168 q169
XSPLIT86 LSmitll_SPLIT 86 q170 q171
XSPLIT87 LSmitll_SPLIT 87 q172 q173
XSPLIT88 LSmitll_SPLIT 88 q174 q175
XSPLIT89 LSmitll_SPLIT 89 q176 q177
XSPLIT90 LSmitll_SPLIT 90 q178 q179
XSPLIT91 LSmitll_SPLIT 91 q180 q181
XSPLIT92 LSmitll_SPLIT 92 q182 q183
XSPLIT93 LSmitll_SPLIT 93 q184 q185
XSPLIT94 LSmitll_SPLIT 94 q186 q187
XSPLIT95 LSmitll_SPLIT 95 q188 q189
XSPLIT96 LSmitll_SPLIT 96 q190 q191
XSPLIT97 LSmitll_SPLIT 97 q192 q193
XSPLIT98 LSmitll_SPLIT 98 q194 q195
XSPLIT99 LSmitll_SPLIT 99 q196 q197
XSPLIT100 LSmitll_SPLIT 100 q198 q199
XSPLIT101 LSmitll_SPLIT 101 q200 q201
XSPLIT102 LSmitll_SPLIT 102 q202 q203
XSPLIT103 LSmitll_SPLIT 103 q204 q205
XSPLIT104 LSmitll_SPLIT 104 q206 q207
XSPLIT105 LSmitll_SPLIT 105 q208 q209
XSPLIT106 LSmitll_SPLIT 106 q210 q211
XSPLIT107 LSmitll_SPLIT 107 q212 q213
XSPLIT108 LSmitll_SPLIT 108 q214 q215
XSPLIT109 LSmitll_SPLIT 109 q216 q217
XSPLIT110 LSmitll_SPLIT 110 q218 q219
XSPLIT111 LSmitll_SPLIT 111 q220 q221
XSPLIT112 LSmitll_SPLIT 112 q222 q223
XSPLIT113 LSmitll_SPLIT 113 q224 q225
XSPLIT114 LSmitll_SPLIT 114 q226 q227
XSPLIT115 LSmitll_SPLIT 115 q228 q229
XSPLIT116 LSmitll_SPLIT 116 q230 q231
XSPLIT117 LSmitll_SPLIT 117 q232 q233
XSPLIT118 LSmitll_SPLIT 118 q234 q235
XSPLIT119 LSmitll_SPLIT 119 q236 q237
XSPLIT120 LSmitll_SPLIT 120 q238 q239
XSPLIT121 LSmitll_SPLIT 121 q240 q241
XSPLIT122 LSmitll_SPLIT 122 q242 q243
XSPLIT123 LSmitll_SPLIT 123 q244 q245
XSPLIT124 LSmitll_SPLIT 124 q246 q247
XSPLIT125 LSmitll_SPLIT 125 q248 q249
XSPLIT126 LSmitll_SPLIT 126 q250 q251
XSPLIT127 LSmitll_SPLIT 127 q252 q253
XSPLIT128 LSmitll_SPLIT 128 q254 q255
XSPLIT129 LSmitll_SPLIT 129 q256 q257
XSPLIT130 LSmitll_SPLIT 130 q258 q259
XSPLIT131 LSmitll_SPLIT 131 q260 q261
XSPLIT132 LSmitll_SPLIT 132 q262 q263
XSPLIT133 LSmitll_SPLIT 133 q264 q265
XSPLIT134 LSmitll_SPLIT 134 q266 q267
XSPLIT135 LSmitll_SPLIT 135 q268 q269
XSPLIT136 LSmitll_SPLIT 136 q270 q271
XSPLIT137 LSmitll_SPLIT 137 q272 q273
XSPLIT138 LSmitll_SPLIT 138 q274 q275
XSPLIT139 LSmitll_SPLIT 139 q276 q277
XSPLIT140 LSmitll_SPLIT 140 q278 q279
XSPLIT141 LSmitll_SPLIT 141 q280 q281
XSPLIT142 LSmitll_SPLIT 142 q282 q283
XSPLIT143 LSmitll_SPLIT 143 q284 q285
XSPLIT144 LSmitll_SPLIT 144 q286 q287
XSPLIT145 LSmitll_SPLIT 145 q288 q289
XSPLIT146 LSmitll_SPLIT 146 q290 q291
XSPLIT147 LSmitll_SPLIT 147 q292 q293
XSPLIT148 LSmitll_SPLIT 148 q294 q295
XSPLIT149 LSmitll_SPLIT 149 q296 q297
XSPLIT150 LSmitll_SPLIT 150 q298 q299
XSPLIT151 LSmitll_SPLIT 151 q300 q301
XSPLIT152 LSmitll_SPLIT 152 q302 q303
XSPLIT153 LSmitll_SPLIT 153 q304 q305
XSPLIT154 LSmitll_SPLIT 154 q306 q307
XSPLIT155 LSmitll_SPLIT 155 q308 q309
XSPLIT156 LSmitll_SPLIT 156 q310 q311
XSPLIT157 LSmitll_SPLIT 157 q312 q313
XSPLIT158 LSmitll_SPLIT 158 q314 q315
XSPLIT159 LSmitll_SPLIT 159 q316 q317
XSPLIT160 LSmitll_SPLIT 160 q318 q319
XSPLIT161 LSmitll_SPLIT 161 q320 q321
XSPLIT162 LSmitll_SPLIT 162 q322 q323
XSPLIT163 LSmitll_SPLIT 163 q324 q325
XSPLIT164 LSmitll_SPLIT 164 q326 q327
XSPLIT165 LSmitll_SPLIT 165 q328 q329
XSPLIT166 LSmitll_SPLIT 166 q330 q331
XSPLIT167 LSmitll_SPLIT 167 q332 q333
XSPLIT168 LSmitll_SPLIT 168 q334 q335
XSPLIT169 LSmitll_SPLIT 169 q336 q337
XSPLIT170 LSmitll_SPLIT 170 q338 q339
XSPLIT171 LSmitll_SPLIT 171 q340 q341
XSPLIT172 LSmitll_SPLIT 172 q342 q343
XSPLIT173 LSmitll_SPLIT 173 q344 q345
XSPLIT174 LSmitll_SPLIT 174 q346 q347
XSPLIT175 LSmitll_SPLIT 175 q348 q349
XSPLIT176 LSmitll_SPLIT 176 q350 q351
XSPLIT177 LSmitll_SPLIT 177 q352 q353
XSPLIT178 LSmitll_SPLIT 178 q354 q355
XSPLIT179 LSmitll_SPLIT 179 q356 q357
XSPLIT180 LSmitll_SPLIT 180 q358 q359
XSPLIT181 LSmitll_SPLIT 181 q360 q361
XSPLIT182 LSmitll_SPLIT 182 q362 q363
XSPLIT183 LSmitll_SPLIT 183 q364 q365
XSPLIT184 LSmitll_SPLIT 184 q366 q367
XSPLIT185 LSmitll_SPLIT 185 q368 q369
XSPLIT186 LSmitll_SPLIT 186 q370 q371
XSPLIT187 LSmitll_SPLIT 187 q372 q373
XSPLIT188 LSmitll_SPLIT 188 q374 q375
XSPLIT189 LSmitll_SPLIT 189 q376 q377
XSPLIT190 LSmitll_SPLIT 190 q378 q379
XSPLIT191 LSmitll_SPLIT 191 q380 q381
XSPLIT192 LSmitll_SPLIT 192 q382 q383
XSPLIT193 LSmitll_SPLIT 193 q384 q385
XSPLIT194 LSmitll_SPLIT 194 q386 q387
XSPLIT195 LSmitll_SPLIT 195 q388 q389
XSPLIT196 LSmitll_SPLIT 196 q390 q391
XSPLIT197 LSmitll_SPLIT 197 q392 q393
XSPLIT198 LSmitll_SPLIT 198 q394 q395
XSPLIT199 LSmitll_SPLIT 199 q396 q397
XSPLIT200 LSmitll_SPLIT 200 q398 q399
XSPLIT201 LSmitll_SPLIT 201 q400 q401
XSPLIT202 LSmitll_SPLIT 202 q402 q403
XSPLIT203 LSmitll_SPLIT 203 q404 q405
XSPLIT204 LSmitll_SPLIT 204 q406 q407
XSPLIT205 LSmitll_SPLIT 205 q408 q409
XSPLIT206 LSmitll_SPLIT 206 q410 q411
XSPLIT207 LSmitll_SPLIT 207 q412 q413
XSPLIT208 LSmitll_SPLIT 208 q414 q415
XSPLIT209 LSmitll_SPLIT 209 q416 q417
XSPLIT210 LSmitll_SPLIT 210 q418 q419
XSPLIT211 LSmitll_SPLIT 211 q420 q421
XSPLIT212 LSmitll_SPLIT 212 q422 q423
XSPLIT213 LSmitll_SPLIT 213 q424 q425
XSPLIT214 LSmitll_SPLIT 214 q426 q427
XSPLIT215 LSmitll_SPLIT 215 q428 q429
XSPLIT216 LSmitll_SPLIT 216 q430 q431
XSPLIT217 LSmitll_SPLIT 217 q432 q433
XSPLIT218 LSmitll_SPLIT 218 q434 q435
XSPLIT219 LSmitll_SPLIT 219 q436 q437
XSPLIT220 LSmitll_SPLIT 220 q438 q439
XSPLIT221 LSmitll_SPLIT 221 q440 q441
XSPLIT222 LSmitll_SPLIT 222 q442 q443
XSPLIT223 LSmitll_SPLIT 223 q444 q445
XSPLIT224 LSmitll_SPLIT 224 q446 q447
XSPLIT225 LSmitll_SPLIT 225 q448 q449
XSPLIT226 LSmitll_SPLIT 226 q450 q451
XSPLIT227 LSmitll_SPLIT 227 q452 q453
XSPLIT228 LSmitll_SPLIT 228 q454 q455
XSPLIT229 LSmitll_SPLIT 229 q456 q457
XSPLIT230 LSmitll_SPLIT 230 q458 q459
XSPLIT231 LSmitll_SPLIT 231 q460 q461
XSPLIT232 LSmitll_SPLIT 232 q462 q463
XSPLIT233 LSmitll_SPLIT 233 q464 q465
XSPLIT234 LSmitll_SPLIT 234 q466 q467
XSPLIT235 LSmitll_SPLIT 235 q468 q469
XSPLIT236 LSmitll_SPLIT 236 q470 q471
XSPLIT237 LSmitll_SPLIT 237 q472 q473
XSPLIT238 LSmitll_SPLIT 238 q474 q475
XSPLIT239 LSmitll_SPLIT 239 q476 q477
XSPLIT240 LSmitll_SPLIT 240 q478 q479
XSPLIT241 LSmitll_SPLIT 241 q480 q481
XSPLIT242 LSmitll_SPLIT 242 q482 q483
XSPLIT243 LSmitll_SPLIT 243 q484 q485
XSPLIT244 LSmitll_SPLIT 244 q486 q487
XSPLIT245 LSmitll_SPLIT 245 q488 q489
XSPLIT246 LSmitll_SPLIT 246 q490 q491
XSPLIT247 LSmitll_SPLIT 247 q492 q493
XSPLIT248 LSmitll_SPLIT 248 q494 q495
XSPLIT249 LSmitll_SPLIT 249 q496 q497
XSPLIT250 LSmitll_SPLIT 250 q498 q499
XSPLIT251 LSmitll_SPLIT 251 q500 q501
XSPLIT252 LSmitll_SPLIT 252 q502 q503
XSPLIT253 LSmitll_SPLIT 253 q504 q505
XSPLIT254 LSmitll_SPLIT 254 q506 q507
XSPLIT255 LSmitll_SPLIT 255 q508 q509
XSPLIT256 LSmitll_SPLIT 256 q510 q511
XSPLIT257 LSmitll_SPLIT 257 q512 q513
XSPLIT258 LSmitll_SPLIT 258 q514 q515
XSPLIT259 LSmitll_SPLIT 259 q516 q517
XSPLIT260 LSmitll_SPLIT 260 q518 q519
XSPLIT261 LSmitll_SPLIT 261 q520 q521
XSPLIT262 LSmitll_SPLIT 262 q522 q523
XSPLIT263 LSmitll_SPLIT 263 q524 q525
XSPLIT264 LSmitll_SPLIT 264 q526 q527
XSPLIT265 LSmitll_SPLIT 265 q528 q529
XSPLIT266 LSmitll_SPLIT 266 q530 q531
XSPLIT267 LSmitll_SPLIT 267 q532 q533
XSPLIT268 LSmitll_SPLIT 268 q534 q535
XSPLIT269 LSmitll_SPLIT 269 q536 q537
XSPLIT270 LSmitll_SPLIT 270 q538 q539
XSPLIT271 LSmitll_SPLIT 271 q540 q541
XSPLIT272 LSmitll_SPLIT 272 q542 q543
XSPLIT273 LSmitll_SPLIT 273 q544 q545
XSPLIT274 LSmitll_SPLIT 274 q546 q547
XSPLIT275 LSmitll_SPLIT 275 q548 q549
XSPLIT276 LSmitll_SPLIT 276 q550 q551
XSPLIT277 LSmitll_SPLIT 277 q552 q553
XSPLIT278 LSmitll_SPLIT 278 q554 q555
XSPLIT279 LSmitll_SPLIT 279 q556 q557
XSPLIT280 LSmitll_SPLIT 280 q558 q559
XSPLIT281 LSmitll_SPLIT 281 q560 q561
XSPLIT282 LSmitll_SPLIT 282 q562 q563
XSPLIT283 LSmitll_SPLIT 283 q564 q565
XSPLIT284 LSmitll_SPLIT 284 q566 q567
XSPLIT285 LSmitll_SPLIT 285 q568 q569
XSPLIT286 LSmitll_SPLIT 286 q570 q571
XSPLIT287 LSmitll_SPLIT 287 q572 q573
XSPLIT288 LSmitll_SPLIT 288 q574 q575
XSPLIT289 LSmitll_SPLIT 289 q576 q577
XSPLIT290 LSmitll_SPLIT 290 q578 q579
XSPLIT291 LSmitll_SPLIT 291 q580 q581
XSPLIT292 LSmitll_SPLIT 292 q582 q583
XSPLIT293 LSmitll_SPLIT 293 q584 q585
XSPLIT294 LSmitll_SPLIT 294 q586 q587
XSPLIT295 LSmitll_SPLIT 295 q588 q589
XSPLIT296 LSmitll_SPLIT 296 q590 q591
XSPLIT297 LSmitll_SPLIT 297 q592 q593
XSPLIT298 LSmitll_SPLIT 298 q594 q595
XSPLIT299 LSmitll_SPLIT 299 q596 q597
XSPLIT300 LSmitll_SPLIT 300 q598 q599
XSPLIT301 LSmitll_SPLIT 301 q600 q601
XSPLIT302 LSmitll_SPLIT 302 q602 q603
XSPLIT303 LSmitll_SPLIT 303 q604 q605
XSPLIT304 LSmitll_SPLIT 304 q606 q607
XSPLIT305 LSmitll_SPLIT 305 q608 q609
XSPLIT306 LSmitll_SPLIT 306 q610 q611
XSPLIT307 LSmitll_SPLIT 307 q612 q613
XSPLIT308 LSmitll_SPLIT 308 q614 q615
XSPLIT309 LSmitll_SPLIT 309 q616 q617
XSPLIT310 LSmitll_SPLIT 310 q618 q619
XSPLIT311 LSmitll_SPLIT 311 q620 q621
XSPLIT312 LSmitll_SPLIT 312 q622 q623
XSPLIT313 LSmitll_SPLIT 313 q624 q625
XSPLIT314 LSmitll_SPLIT 314 q626 q627
XSPLIT315 LSmitll_SPLIT 315 q628 q629
XSPLIT316 LSmitll_SPLIT 316 q630 q631
XSPLIT317 LSmitll_SPLIT 317 q632 q633
XSPLIT318 LSmitll_SPLIT 318 q634 q635
XSPLIT319 LSmitll_SPLIT 319 q636 q637
XSPLIT320 LSmitll_SPLIT 320 q638 q639
XSPLIT321 LSmitll_SPLIT 321 q640 q641
XSPLIT322 LSmitll_SPLIT 322 q642 q643
XSPLIT323 LSmitll_SPLIT 323 q644 q645
XSPLIT324 LSmitll_SPLIT 324 q646 q647
XSPLIT325 LSmitll_SPLIT 325 q648 q649
XSPLIT326 LSmitll_SPLIT 326 q650 q651
XSPLIT327 LSmitll_SPLIT 327 q652 q653
XSPLIT328 LSmitll_SPLIT 328 q654 q655
XSPLIT329 LSmitll_SPLIT 329 q656 q657
XSPLIT330 LSmitll_SPLIT 330 q658 q659
XSPLIT331 LSmitll_SPLIT 331 q660 q661
XSPLIT332 LSmitll_SPLIT 332 q662 q663
XSPLIT333 LSmitll_SPLIT 333 q664 q665
XSPLIT334 LSmitll_SPLIT 334 q666 q667
XSPLIT335 LSmitll_SPLIT 335 q668 q669
XSPLIT336 LSmitll_SPLIT 336 q670 q671
XSPLIT337 LSmitll_SPLIT 337 q672 q673
XSPLIT338 LSmitll_SPLIT 338 q674 q675
XSPLIT339 LSmitll_SPLIT 339 q676 q677
XSPLIT340 LSmitll_SPLIT 340 q678 q679
XSPLIT341 LSmitll_SPLIT 341 q680 q681
XSPLIT342 LSmitll_SPLIT 342 q682 q683
XSPLIT343 LSmitll_SPLIT 343 q684 q685
XSPLIT344 LSmitll_SPLIT 344 q686 q687
XSPLIT345 LSmitll_SPLIT 345 q688 q689
XSPLIT346 LSmitll_SPLIT 346 q690 q691
XSPLIT347 LSmitll_SPLIT 347 q692 q693
XSPLIT348 LSmitll_SPLIT 348 q694 q695
XSPLIT349 LSmitll_SPLIT 349 q696 q697
XSPLIT350 LSmitll_SPLIT 350 q698 q699
XSPLIT351 LSmitll_SPLIT 351 q700 q701
XSPLIT352 LSmitll_SPLIT 352 q702 q703
XSPLIT353 LSmitll_SPLIT 353 q704 q705
XSPLIT354 LSmitll_SPLIT 354 q706 q707
XSPLIT355 LSmitll_SPLIT 355 q708 q709
XSPLIT356 LSmitll_SPLIT 356 q710 q711
XSPLIT357 LSmitll_SPLIT 357 q712 q713
XSPLIT358 LSmitll_SPLIT 358 q714 q715
XSPLIT359 LSmitll_SPLIT 359 q716 q717
XSPLIT360 LSmitll_SPLIT 360 q718 q719
XSPLIT361 LSmitll_SPLIT 361 q720 q721
XSPLIT362 LSmitll_SPLIT 362 q722 q723
XSPLIT363 LSmitll_SPLIT 363 q724 q725
XSPLIT364 LSmitll_SPLIT 364 q726 q727
XSPLIT365 LSmitll_SPLIT 365 q728 q729
XSPLIT366 LSmitll_SPLIT 366 q730 q731
XSPLIT367 LSmitll_SPLIT 367 q732 q733
XSPLIT368 LSmitll_SPLIT 368 q734 q735
XSPLIT369 LSmitll_SPLIT 369 q736 q737
XSPLIT370 LSmitll_SPLIT 370 q738 q739
XSPLIT371 LSmitll_SPLIT 371 q740 q741
XSPLIT372 LSmitll_SPLIT 372 q742 q743
XSPLIT373 LSmitll_SPLIT 373 q744 q745
XSPLIT374 LSmitll_SPLIT 374 q746 q747
XSPLIT375 LSmitll_SPLIT 375 q748 q749
XSPLIT376 LSmitll_SPLIT 376 q750 q751
XSPLIT377 LSmitll_SPLIT 377 q752 q753
XSPLIT378 LSmitll_SPLIT 378 q754 q755
XSPLIT379 LSmitll_SPLIT 379 q756 q757
XSPLIT380 LSmitll_SPLIT 380 q758 q759
XSPLIT381 LSmitll_SPLIT 381 q760 q761
XSPLIT382 LSmitll_SPLIT 382 q762 q763
XSPLIT383 LSmitll_SPLIT 383 q764 q765
XSPLIT384 LSmitll_SPLIT 384 q766 q767
XSPLIT385 LSmitll_SPLIT 385 q768 q769
XSPLIT386 LSmitll_SPLIT 386 q770 q771
XSPLIT387 LSmitll_SPLIT 387 q772 q773
XSPLIT388 LSmitll_SPLIT 388 q774 q775
XSPLIT389 LSmitll_SPLIT 389 q776 q777
XSPLIT390 LSmitll_SPLIT 390 q778 q779
XSPLIT391 LSmitll_SPLIT 391 q780 q781
XSPLIT392 LSmitll_SPLIT 392 q782 q783
XSPLIT393 LSmitll_SPLIT 393 q784 q785
XSPLIT394 LSmitll_SPLIT 394 q786 q787
XSPLIT395 LSmitll_SPLIT 395 q788 q789
XSPLIT396 LSmitll_SPLIT 396 q790 q791
XSPLIT397 LSmitll_SPLIT 397 q792 q793
XSPLIT398 LSmitll_SPLIT 398 q794 q795
XSPLIT399 LSmitll_SPLIT 399 q796 q797
XSPLIT400 LSmitll_SPLIT 400 q798 q799
XSPLIT401 LSmitll_SPLIT 401 q800 q801
XSPLIT402 LSmitll_SPLIT 402 q802 q803
XSPLIT403 LSmitll_SPLIT 403 q804 q805
XSPLIT404 LSmitll_SPLIT 404 q806 q807
XSPLIT405 LSmitll_SPLIT 405 q808 q809
XSPLIT406 LSmitll_SPLIT 406 q810 q811
XSPLIT407 LSmitll_SPLIT 407 q812 q813
XSPLIT408 LSmitll_SPLIT 408 q814 q815
XSPLIT409 LSmitll_SPLIT 409 q816 q817
XSPLIT410 LSmitll_SPLIT 410 q818 q819
XSPLIT411 LSmitll_SPLIT 411 q820 q821
XSPLIT412 LSmitll_SPLIT 412 q822 q823
XSPLIT413 LSmitll_SPLIT 413 q824 q825
XSPLIT414 LSmitll_SPLIT 414 q826 q827
XSPLIT415 LSmitll_SPLIT 415 q828 q829
XSPLIT416 LSmitll_SPLIT 416 q830 q831
XSPLIT417 LSmitll_SPLIT 417 q832 q833
XSPLIT418 LSmitll_SPLIT 418 q834 q835
XSPLIT419 LSmitll_SPLIT 419 q836 q837
XSPLIT420 LSmitll_SPLIT 420 q838 q839
XSPLIT421 LSmitll_SPLIT 421 q840 q841
XSPLIT422 LSmitll_SPLIT 422 q842 q843
XSPLIT423 LSmitll_SPLIT 423 q844 q845
XSPLIT424 LSmitll_SPLIT 424 q846 q847
XSPLIT425 LSmitll_SPLIT 425 q848 q849
XSPLIT426 LSmitll_SPLIT 426 q850 q851
XSPLIT427 LSmitll_SPLIT 427 q852 q853
XSPLIT428 LSmitll_SPLIT 428 q854 q855
XSPLIT429 LSmitll_SPLIT 429 q856 q857
XSPLIT430 LSmitll_SPLIT 430 q858 q859
XSPLIT431 LSmitll_SPLIT 431 q860 q861
XSPLIT432 LSmitll_SPLIT 432 q862 q863
XSPLIT433 LSmitll_SPLIT 433 q864 q865
XSPLIT434 LSmitll_SPLIT 434 q866 q867
XSPLIT435 LSmitll_SPLIT 435 q868 q869
XSPLIT436 LSmitll_SPLIT 436 q870 q871
XSPLIT437 LSmitll_SPLIT 437 q872 q873
XSPLIT438 LSmitll_SPLIT 438 q874 q875
XSPLIT439 LSmitll_SPLIT 439 q876 q877
XSPLIT440 LSmitll_SPLIT 440 q878 q879
XSPLIT441 LSmitll_SPLIT 441 q880 q881
XSPLIT442 LSmitll_SPLIT 442 q882 q883
XSPLIT443 LSmitll_SPLIT 443 q884 q885
XSPLIT444 LSmitll_SPLIT 444 q886 q887
XSPLIT445 LSmitll_SPLIT 445 q888 q889
XSPLIT446 LSmitll_SPLIT 446 q890 q891
XSPLIT447 LSmitll_SPLIT 447 q892 q893
XSPLIT448 LSmitll_SPLIT 448 q894 q895
XSPLIT449 LSmitll_SPLIT 449 q896 q897
XSPLIT450 LSmitll_SPLIT 450 q898 q899
XSPLIT451 LSmitll_SPLIT 451 q900 q901
XSPLIT452 LSmitll_SPLIT 452 q902 q903
XSPLIT453 LSmitll_SPLIT 453 q904 q905
XSPLIT454 LSmitll_SPLIT 454 q906 q907
XSPLIT455 LSmitll_SPLIT 455 q908 q909
XSPLIT456 LSmitll_SPLIT 456 q910 q911
XSPLIT457 LSmitll_SPLIT 457 q912 q913
XSPLIT458 LSmitll_SPLIT 458 q914 q915
XSPLIT459 LSmitll_SPLIT 459 q916 q917
XSPLIT460 LSmitll_SPLIT 460 q918 q919
XSPLIT461 LSmitll_SPLIT 461 q920 q921
XSPLIT462 LSmitll_SPLIT 462 q922 q923
XSPLIT463 LSmitll_SPLIT 463 q924 q925
XSPLIT464 LSmitll_SPLIT 464 q926 q927
XSPLIT465 LSmitll_SPLIT 465 q928 q929
XSPLIT466 LSmitll_SPLIT 466 q930 q931
XSPLIT467 LSmitll_SPLIT 467 q932 q933
XSPLIT468 LSmitll_SPLIT 468 q934 q935
XSPLIT469 LSmitll_SPLIT 469 q936 q937
XSPLIT470 LSmitll_SPLIT 470 q938 q939
XSPLIT471 LSmitll_SPLIT 471 q940 q941
XSPLIT472 LSmitll_SPLIT 472 q942 q943
XSPLIT473 LSmitll_SPLIT 473 q944 q945
XSPLIT474 LSmitll_SPLIT 474 q946 q947
XSPLIT475 LSmitll_SPLIT 475 q948 q949
XSPLIT476 LSmitll_SPLIT 476 q950 q951
XSPLIT477 LSmitll_SPLIT 477 q952 q953
XSPLIT478 LSmitll_SPLIT 478 q954 q955
XSPLIT479 LSmitll_SPLIT 479 q956 q957
XSPLIT480 LSmitll_SPLIT 480 q958 q959
XSPLIT481 LSmitll_SPLIT 481 q960 q961
XSPLIT482 LSmitll_SPLIT 482 q962 q963
XSPLIT483 LSmitll_SPLIT 483 q964 q965
XSPLIT484 LSmitll_SPLIT 484 q966 q967
XSPLIT485 LSmitll_SPLIT 485 q968 q969
XSPLIT486 LSmitll_SPLIT 486 q970 q971
XSPLIT487 LSmitll_SPLIT 487 q972 q973
XSPLIT488 LSmitll_SPLIT 488 q974 q975
XSPLIT489 LSmitll_SPLIT 489 q976 q977
XSPLIT490 LSmitll_SPLIT 490 q978 q979
XSPLIT491 LSmitll_SPLIT 491 q980 q981
XSPLIT492 LSmitll_SPLIT 492 q982 q983
XSPLIT493 LSmitll_SPLIT 493 q984 q985
XSPLIT494 LSmitll_SPLIT 494 q986 q987
XSPLIT495 LSmitll_SPLIT 495 q988 q989
XSPLIT496 LSmitll_SPLIT 496 q990 q991
XSPLIT497 LSmitll_SPLIT 497 q992 q993
XSPLIT498 LSmitll_SPLIT 498 q994 q995
XSPLIT499 LSmitll_SPLIT 499 q996 q997
XSPLIT500 LSmitll_SPLIT 500 q998 q999
XSPLIT501 LSmitll_SPLIT 501 q1000 q1001
XSPLIT502 LSmitll_SPLIT 502 q1002 q1003
XSPLIT503 LSmitll_SPLIT 503 q1004 q1005
XSPLIT504 LSmitll_SPLIT 504 q1006 q1007
XSPLIT505 LSmitll_SPLIT 505 q1008 q1009
XSPLIT506 LSmitll_SPLIT 506 q1010 q1011
XSPLIT507 LSmitll_SPLIT 507 q1012 q1013
XSPLIT508 LSmitll_SPLIT 508 q1014 q1015
XSPLIT509 LSmitll_SPLIT 509 q1016 q1017
XSPLIT510 LSmitll_SPLIT 510 q1018 q1019
XSPLIT511 LSmitll_SPLIT 511 q1020 q1021
XSPLIT512 LSmitll_SPLIT 512 q1022 q1023
XSPLIT513 LSmitll_SPLIT 513 q1024 q1025
XSPLIT514 LSmitll_SPLIT 514 q1026 q1027
XSPLIT515 LSmitll_SPLIT 515 q1028 q1029
XSPLIT516 LSmitll_SPLIT 516 q1030 q1031
XSPLIT517 LSmitll_SPLIT 517 q1032 q1033
XSPLIT518 LSmitll_SPLIT 518 q1034 q1035
XSPLIT519 LSmitll_SPLIT 519 q1036 q1037
XSPLIT520 LSmitll_SPLIT 520 q1038 q1039
XSPLIT521 LSmitll_SPLIT 521 q1040 q1041
XSPLIT522 LSmitll_SPLIT 522 q1042 q1043
XSPLIT523 LSmitll_SPLIT 523 q1044 q1045
XSPLIT524 LSmitll_SPLIT 524 q1046 q1047
XSPLIT525 LSmitll_SPLIT 525 q1048 q1049
XSPLIT526 LSmitll_SPLIT 526 q1050 q1051
XSPLIT527 LSmitll_SPLIT 527 q1052 q1053
XSPLIT528 LSmitll_SPLIT 528 q1054 q1055
XSPLIT529 LSmitll_SPLIT 529 q1056 q1057
XSPLIT530 LSmitll_SPLIT 530 q1058 q1059
XSPLIT531 LSmitll_SPLIT 531 q1060 q1061
XSPLIT532 LSmitll_SPLIT 532 q1062 q1063
XSPLIT533 LSmitll_SPLIT 533 q1064 q1065
XSPLIT534 LSmitll_SPLIT 534 q1066 q1067
XSPLIT535 LSmitll_SPLIT 535 q1068 q1069
XSPLIT536 LSmitll_SPLIT 536 q1070 q1071
XSPLIT537 LSmitll_SPLIT 537 q1072 q1073
XSPLIT538 LSmitll_SPLIT 538 q1074 q1075
XSPLIT539 LSmitll_SPLIT 539 q1076 q1077
XSPLIT540 LSmitll_SPLIT 540 q1078 q1079
XSPLIT541 LSmitll_SPLIT 541 q1080 q1081
XSPLIT542 LSmitll_SPLIT 542 q1082 q1083
XSPLIT543 LSmitll_SPLIT 543 q1084 q1085
XSPLIT544 LSmitll_SPLIT 544 q1086 q1087
XSPLIT545 LSmitll_SPLIT 545 q1088 q1089
XSPLIT546 LSmitll_SPLIT 546 q1090 q1091
XSPLIT547 LSmitll_SPLIT 547 q1092 q1093
XSPLIT548 LSmitll_SPLIT 548 q1094 q1095
XSPLIT549 LSmitll_SPLIT 549 q1096 q1097
XSPLIT550 LSmitll_SPLIT 550 q1098 q1099
XSPLIT551 LSmitll_SPLIT 551 q1100 q1101
XSPLIT552 LSmitll_SPLIT 552 q1102 q1103
XSPLIT553 LSmitll_SPLIT 553 q1104 q1105
XSPLIT554 LSmitll_SPLIT 554 q1106 q1107
XSPLIT555 LSmitll_SPLIT 555 q1108 q1109
XSPLIT556 LSmitll_SPLIT 556 q1110 q1111
XSPLIT557 LSmitll_SPLIT 557 q1112 q1113
XSPLIT558 LSmitll_SPLIT 558 q1114 q1115
XSPLIT559 LSmitll_SPLIT 559 q1116 q1117
XSPLIT560 LSmitll_SPLIT 560 q1118 q1119
XSPLIT561 LSmitll_SPLIT 561 q1120 q1121
XSPLIT562 LSmitll_SPLIT 562 q1122 q1123
XSPLIT563 LSmitll_SPLIT 563 q1124 q1125
XSPLIT564 LSmitll_SPLIT 564 q1126 q1127
XSPLIT565 LSmitll_SPLIT 565 q1128 q1129
XSPLIT566 LSmitll_SPLIT 566 q1130 q1131
XSPLIT567 LSmitll_SPLIT 567 q1132 q1133
XSPLIT568 LSmitll_SPLIT 568 q1134 q1135
XSPLIT569 LSmitll_SPLIT 569 q1136 q1137
XSPLIT570 LSmitll_SPLIT 570 q1138 q1139
XSPLIT571 LSmitll_SPLIT 571 q1140 q1141
XSPLIT572 LSmitll_SPLIT 572 q1142 q1143
XSPLIT573 LSmitll_SPLIT 573 q1144 q1145
XSPLIT574 LSmitll_SPLIT 574 q1146 q1147
XSPLIT575 LSmitll_SPLIT 575 q1148 q1149
XSPLIT576 LSmitll_SPLIT 576 q1150 q1151
XSPLIT577 LSmitll_SPLIT 577 q1152 q1153
XSPLIT578 LSmitll_SPLIT 578 q1154 q1155
XSPLIT579 LSmitll_SPLIT 579 q1156 q1157
XSPLIT580 LSmitll_SPLIT 580 q1158 q1159
XSPLIT581 LSmitll_SPLIT 581 q1160 q1161
XSPLIT582 LSmitll_SPLIT 582 q1162 q1163
XSPLIT583 LSmitll_SPLIT 583 q1164 q1165
XSPLIT584 LSmitll_SPLIT 584 q1166 q1167
XSPLIT585 LSmitll_SPLIT 585 q1168 q1169
XSPLIT586 LSmitll_SPLIT 586 q1170 q1171
XSPLIT587 LSmitll_SPLIT 587 q1172 q1173
XSPLIT588 LSmitll_SPLIT 588 q1174 q1175
XSPLIT589 LSmitll_SPLIT 589 q1176 q1177
XSPLIT590 LSmitll_SPLIT 590 q1178 q1179
XSPLIT591 LSmitll_SPLIT 591 q1180 q1181
XSPLIT592 LSmitll_SPLIT 592 q1182 q1183
XSPLIT593 LSmitll_SPLIT 593 q1184 q1185
XSPLIT594 LSmitll_SPLIT 594 q1186 q1187
XSPLIT595 LSmitll_SPLIT 595 q1188 q1189
XSPLIT596 LSmitll_SPLIT 596 q1190 q1191
XSPLIT597 LSmitll_SPLIT 597 q1192 q1193
XSPLIT598 LSmitll_SPLIT 598 q1194 q1195
XSPLIT599 LSmitll_SPLIT 599 q1196 q1197
XSPLIT600 LSmitll_SPLIT 600 q1198 q1199
XSPLIT601 LSmitll_SPLIT 601 q1200 q1201
XSPLIT602 LSmitll_SPLIT 602 q1202 q1203
XSPLIT603 LSmitll_SPLIT 603 q1204 q1205
XSPLIT604 LSmitll_SPLIT 604 q1206 q1207
XSPLIT605 LSmitll_SPLIT 605 q1208 q1209
XSPLIT606 LSmitll_SPLIT 606 q1210 q1211
XSPLIT607 LSmitll_SPLIT 607 q1212 q1213
XSPLIT608 LSmitll_SPLIT 608 q1214 q1215
XSPLIT609 LSmitll_SPLIT 609 q1216 q1217
XSPLIT610 LSmitll_SPLIT 610 q1218 q1219
XSPLIT611 LSmitll_SPLIT 611 q1220 q1221
XSPLIT612 LSmitll_SPLIT 612 q1222 q1223
XSPLIT613 LSmitll_SPLIT 613 q1224 q1225
XSPLIT614 LSmitll_SPLIT 614 q1226 q1227
XSPLIT615 LSmitll_SPLIT 615 q1228 q1229
XSPLIT616 LSmitll_SPLIT 616 q1230 q1231
XSPLIT617 LSmitll_SPLIT 617 q1232 q1233
XSPLIT618 LSmitll_SPLIT 618 q1234 q1235
XSPLIT619 LSmitll_SPLIT 619 q1236 q1237
XSPLIT620 LSmitll_SPLIT 620 q1238 q1239
XSPLIT621 LSmitll_SPLIT 621 q1240 q1241
XSPLIT622 LSmitll_SPLIT 622 q1242 q1243
XSPLIT623 LSmitll_SPLIT 623 q1244 q1245
XSPLIT624 LSmitll_SPLIT 624 q1246 q1247
XSPLIT625 LSmitll_SPLIT 625 q1248 q1249
XSPLIT626 LSmitll_SPLIT 626 q1250 q1251
XSPLIT627 LSmitll_SPLIT 627 q1252 q1253
XSPLIT628 LSmitll_SPLIT 628 q1254 q1255
XSPLIT629 LSmitll_SPLIT 629 q1256 q1257
XSPLIT630 LSmitll_SPLIT 630 q1258 q1259
XSPLIT631 LSmitll_SPLIT 631 q1260 q1261
XSPLIT632 LSmitll_SPLIT 632 q1262 q1263
XSPLIT633 LSmitll_SPLIT 633 q1264 q1265
XSPLIT634 LSmitll_SPLIT 634 q1266 q1267
XSPLIT635 LSmitll_SPLIT 635 q1268 q1269
XSPLIT636 LSmitll_SPLIT 636 q1270 q1271
XSPLIT637 LSmitll_SPLIT 637 q1272 q1273
XSPLIT638 LSmitll_SPLIT 638 q1274 q1275
XSPLIT639 LSmitll_SPLIT 639 q1276 q1277
XSPLIT640 LSmitll_SPLIT 640 q1278 q1279
XSPLIT641 LSmitll_SPLIT 641 q1280 q1281
XSPLIT642 LSmitll_SPLIT 642 q1282 q1283
XSPLIT643 LSmitll_SPLIT 643 q1284 q1285
XSPLIT644 LSmitll_SPLIT 644 q1286 q1287
XSPLIT645 LSmitll_SPLIT 645 q1288 q1289
XSPLIT646 LSmitll_SPLIT 646 q1290 q1291
XSPLIT647 LSmitll_SPLIT 647 q1292 q1293
XSPLIT648 LSmitll_SPLIT 648 q1294 q1295
XSPLIT649 LSmitll_SPLIT 649 q1296 q1297
XSPLIT650 LSmitll_SPLIT 650 q1298 q1299
XSPLIT651 LSmitll_SPLIT 651 q1300 q1301
XSPLIT652 LSmitll_SPLIT 652 q1302 q1303
XSPLIT653 LSmitll_SPLIT 653 q1304 q1305
XSPLIT654 LSmitll_SPLIT 654 q1306 q1307
XSPLIT655 LSmitll_SPLIT 655 q1308 q1309
XSPLIT656 LSmitll_SPLIT 656 q1310 q1311
XSPLIT657 LSmitll_SPLIT 657 q1312 q1313
XSPLIT658 LSmitll_SPLIT 658 q1314 q1315
XSPLIT659 LSmitll_SPLIT 659 q1316 q1317
XSPLIT660 LSmitll_SPLIT 660 q1318 q1319
XSPLIT661 LSmitll_SPLIT 661 q1320 q1321
XSPLIT662 LSmitll_SPLIT 662 q1322 q1323
XSPLIT663 LSmitll_SPLIT 663 q1324 q1325
XSPLIT664 LSmitll_SPLIT 664 q1326 q1327
XSPLIT665 LSmitll_SPLIT 665 q1328 q1329
XSPLIT666 LSmitll_SPLIT 666 q1330 q1331
XSPLIT667 LSmitll_SPLIT 667 q1332 q1333
XSPLIT668 LSmitll_SPLIT 668 q1334 q1335
XSPLIT669 LSmitll_SPLIT 669 q1336 q1337
XSPLIT670 LSmitll_SPLIT 670 q1338 q1339
XSPLIT671 LSmitll_SPLIT 671 q1340 q1341
XSPLIT672 LSmitll_SPLIT 672 q1342 q1343
XSPLIT673 LSmitll_SPLIT 673 q1344 q1345
XSPLIT674 LSmitll_SPLIT 674 q1346 q1347
XSPLIT675 LSmitll_SPLIT 675 q1348 q1349
XSPLIT676 LSmitll_SPLIT 676 q1350 q1351
XSPLIT677 LSmitll_SPLIT 677 q1352 q1353
XSPLIT678 LSmitll_SPLIT 678 q1354 q1355
XSPLIT679 LSmitll_SPLIT 679 q1356 q1357
XSPLIT680 LSmitll_SPLIT 680 q1358 q1359
XSPLIT681 LSmitll_SPLIT 681 q1360 q1361
XSPLIT682 LSmitll_SPLIT 682 q1362 q1363
XSPLIT683 LSmitll_SPLIT 683 q1364 q1365
XSPLIT684 LSmitll_SPLIT 684 q1366 q1367
XSPLIT685 LSmitll_SPLIT 685 q1368 q1369
XSPLIT686 LSmitll_SPLIT 686 q1370 q1371
XSPLIT687 LSmitll_SPLIT 687 q1372 q1373
XSPLIT688 LSmitll_SPLIT 688 q1374 q1375
XSPLIT689 LSmitll_SPLIT 689 q1376 q1377
XSPLIT690 LSmitll_SPLIT 690 q1378 q1379
XSPLIT691 LSmitll_SPLIT 691 q1380 q1381
XSPLIT692 LSmitll_SPLIT 692 q1382 q1383
XSPLIT693 LSmitll_SPLIT 693 q1384 q1385
XSPLIT694 LSmitll_SPLIT 694 q1386 q1387
XSPLIT695 LSmitll_SPLIT 695 q1388 q1389
XSPLIT696 LSmitll_SPLIT 696 q1390 q1391
XSPLIT697 LSmitll_SPLIT 697 q1392 q1393
XSPLIT698 LSmitll_SPLIT 698 q1394 q1395
XSPLIT699 LSmitll_SPLIT 699 q1396 q1397
XSPLIT700 LSmitll_SPLIT 700 q1398 q1399
XSPLIT701 LSmitll_SPLIT 701 q1400 q1401
XSPLIT702 LSmitll_SPLIT 702 q1402 q1403
XSPLIT703 LSmitll_SPLIT 703 q1404 q1405
XSPLIT704 LSmitll_SPLIT 704 q1406 q1407
XSPLIT705 LSmitll_SPLIT 705 q1408 q1409
XSPLIT706 LSmitll_SPLIT 706 q1410 q1411
XSPLIT707 LSmitll_SPLIT 707 q1412 q1413
XSPLIT708 LSmitll_SPLIT 708 q1414 q1415
XSPLIT709 LSmitll_SPLIT 709 q1416 q1417
XSPLIT710 LSmitll_SPLIT 710 q1418 q1419
XSPLIT711 LSmitll_SPLIT 711 q1420 q1421
XSPLIT712 LSmitll_SPLIT 712 q1422 q1423
XSPLIT713 LSmitll_SPLIT 713 q1424 q1425
XSPLIT714 LSmitll_SPLIT 714 q1426 q1427
XSPLIT715 LSmitll_SPLIT 715 q1428 q1429
XSPLIT716 LSmitll_SPLIT 716 q1430 q1431
XSPLIT717 LSmitll_SPLIT 717 q1432 q1433
XSPLIT718 LSmitll_SPLIT 718 q1434 q1435
XSPLIT719 LSmitll_SPLIT 719 q1436 q1437
XSPLIT720 LSmitll_SPLIT 720 q1438 q1439
XSPLIT721 LSmitll_SPLIT 721 q1440 q1441
XSPLIT722 LSmitll_SPLIT 722 q1442 q1443
XSPLIT723 LSmitll_SPLIT 723 q1444 q1445
XSPLIT724 LSmitll_SPLIT 724 q1446 q1447
XSPLIT725 LSmitll_SPLIT 725 q1448 q1449
XSPLIT726 LSmitll_SPLIT 726 q1450 q1451
XSPLIT727 LSmitll_SPLIT 727 q1452 q1453
XSPLIT728 LSmitll_SPLIT 728 q1454 q1455
XSPLIT729 LSmitll_SPLIT 729 q1456 q1457
XSPLIT730 LSmitll_SPLIT 730 q1458 q1459
XSPLIT731 LSmitll_SPLIT 731 q1460 q1461
XSPLIT732 LSmitll_SPLIT 732 q1462 q1463
XSPLIT733 LSmitll_SPLIT 733 q1464 q1465
XSPLIT734 LSmitll_SPLIT 734 q1466 q1467
XSPLIT735 LSmitll_SPLIT 735 q1468 q1469
XSPLIT736 LSmitll_SPLIT 736 q1470 q1471
XSPLIT737 LSmitll_SPLIT 737 q1472 q1473
XSPLIT738 LSmitll_SPLIT 738 q1474 q1475
XSPLIT739 LSmitll_SPLIT 739 q1476 q1477
XSPLIT740 LSmitll_SPLIT 740 q1478 q1479
XSPLIT741 LSmitll_SPLIT 741 q1480 q1481
XSPLIT742 LSmitll_SPLIT 742 q1482 q1483
XSPLIT743 LSmitll_SPLIT 743 q1484 q1485
XSPLIT744 LSmitll_SPLIT 744 q1486 q1487
XSPLIT745 LSmitll_SPLIT 745 q1488 q1489
XSPLIT746 LSmitll_SPLIT 746 q1490 q1491
XSPLIT747 LSmitll_SPLIT 747 q1492 q1493
XSPLIT748 LSmitll_SPLIT 748 q1494 q1495
XSPLIT749 LSmitll_SPLIT 749 q1496 q1497
XSPLIT750 LSmitll_SPLIT 750 q1498 q1499
XSPLIT751 LSmitll_SPLIT 751 q1500 q1501
XSPLIT752 LSmitll_SPLIT 752 q1502 q1503
XSPLIT753 LSmitll_SPLIT 753 q1504 q1505
XSPLIT754 LSmitll_SPLIT 754 q1506 q1507
XSPLIT755 LSmitll_SPLIT 755 q1508 q1509
XSPLIT756 LSmitll_SPLIT 756 q1510 q1511
XSPLIT757 LSmitll_SPLIT 757 q1512 q1513
XSPLIT758 LSmitll_SPLIT 758 q1514 q1515
XSPLIT759 LSmitll_SPLIT 759 q1516 q1517
XSPLIT760 LSmitll_SPLIT 760 q1518 q1519
XSPLIT761 LSmitll_SPLIT 761 q1520 q1521
XSPLIT762 LSmitll_SPLIT 762 q1522 q1523
XSPLIT763 LSmitll_SPLIT 763 q1524 q1525
XSPLIT764 LSmitll_SPLIT 764 q1526 q1527
XSPLIT765 LSmitll_SPLIT 765 q1528 q1529
XSPLIT766 LSmitll_SPLIT 766 q1530 q1531
XSPLIT767 LSmitll_SPLIT 767 q1532 q1533
XSPLIT768 LSmitll_SPLIT 768 q1534 q1535
XSPLIT769 LSmitll_SPLIT 769 q1536 q1537
XSPLIT770 LSmitll_SPLIT 770 q1538 q1539
XSPLIT771 LSmitll_SPLIT 771 q1540 q1541
XSPLIT772 LSmitll_SPLIT 772 q1542 q1543
XSPLIT773 LSmitll_SPLIT 773 q1544 q1545
XSPLIT774 LSmitll_SPLIT 774 q1546 q1547
XSPLIT775 LSmitll_SPLIT 775 q1548 q1549
XSPLIT776 LSmitll_SPLIT 776 q1550 q1551
XSPLIT777 LSmitll_SPLIT 777 q1552 q1553
XSPLIT778 LSmitll_SPLIT 778 q1554 q1555
XSPLIT779 LSmitll_SPLIT 779 q1556 q1557
XSPLIT780 LSmitll_SPLIT 780 q1558 q1559
XSPLIT781 LSmitll_SPLIT 781 q1560 q1561
XSPLIT782 LSmitll_SPLIT 782 q1562 q1563
XSPLIT783 LSmitll_SPLIT 783 q1564 q1565
XSPLIT784 LSmitll_SPLIT 784 q1566 q1567
XSPLIT785 LSmitll_SPLIT 785 q1568 q1569
XSPLIT786 LSmitll_SPLIT 786 q1570 q1571
XSPLIT787 LSmitll_SPLIT 787 q1572 q1573
XSPLIT788 LSmitll_SPLIT 788 q1574 q1575
XSPLIT789 LSmitll_SPLIT 789 q1576 q1577
XSPLIT790 LSmitll_SPLIT 790 q1578 q1579
XSPLIT791 LSmitll_SPLIT 791 q1580 q1581
XSPLIT792 LSmitll_SPLIT 792 q1582 q1583
XSPLIT793 LSmitll_SPLIT 793 q1584 q1585
XSPLIT794 LSmitll_SPLIT 794 q1586 q1587
XSPLIT795 LSmitll_SPLIT 795 q1588 q1589
XSPLIT796 LSmitll_SPLIT 796 q1590 q1591
XSPLIT797 LSmitll_SPLIT 797 q1592 q1593
XSPLIT798 LSmitll_SPLIT 798 q1594 q1595
XSPLIT799 LSmitll_SPLIT 799 q1596 q1597
XSPLIT800 LSmitll_SPLIT 800 q1598 q1599
XSPLIT801 LSmitll_SPLIT 801 q1600 q1601
XSPLIT802 LSmitll_SPLIT 802 q1602 q1603
XSPLIT803 LSmitll_SPLIT 803 q1604 q1605
XSPLIT804 LSmitll_SPLIT 804 q1606 q1607
XSPLIT805 LSmitll_SPLIT 805 q1608 q1609
XSPLIT806 LSmitll_SPLIT 806 q1610 q1611
XSPLIT807 LSmitll_SPLIT 807 q1612 q1613
XSPLIT808 LSmitll_SPLIT 808 q1614 q1615
XSPLIT809 LSmitll_SPLIT 809 q1616 q1617
XSPLIT810 LSmitll_SPLIT 810 q1618 q1619
XSPLIT811 LSmitll_SPLIT 811 q1620 q1621
XSPLIT812 LSmitll_SPLIT 812 q1622 q1623
XSPLIT813 LSmitll_SPLIT 813 q1624 q1625
XSPLIT814 LSmitll_SPLIT 814 q1626 q1627
XSPLIT815 LSmitll_SPLIT 815 q1628 q1629
XSPLIT816 LSmitll_SPLIT 816 q1630 q1631
XSPLIT817 LSmitll_SPLIT 817 q1632 q1633
XSPLIT818 LSmitll_SPLIT 818 q1634 q1635
XSPLIT819 LSmitll_SPLIT 819 q1636 q1637
XSPLIT820 LSmitll_SPLIT 820 q1638 q1639
XSPLIT821 LSmitll_SPLIT 821 q1640 q1641
XSPLIT822 LSmitll_SPLIT 822 q1642 q1643
XSPLIT823 LSmitll_SPLIT 823 q1644 q1645
XSPLIT824 LSmitll_SPLIT 824 q1646 q1647
XSPLIT825 LSmitll_SPLIT 825 q1648 q1649
XSPLIT826 LSmitll_SPLIT 826 q1650 q1651
XSPLIT827 LSmitll_SPLIT 827 q1652 q1653
XSPLIT828 LSmitll_SPLIT 828 q1654 q1655
XSPLIT829 LSmitll_SPLIT 829 q1656 q1657
XSPLIT830 LSmitll_SPLIT 830 q1658 q1659
XSPLIT831 LSmitll_SPLIT 831 q1660 q1661
XSPLIT832 LSmitll_SPLIT 832 q1662 q1663
XSPLIT833 LSmitll_SPLIT 833 q1664 q1665
XSPLIT834 LSmitll_SPLIT 834 q1666 q1667
XSPLIT835 LSmitll_SPLIT 835 q1668 q1669
XSPLIT836 LSmitll_SPLIT 836 q1670 q1671
XSPLIT837 LSmitll_SPLIT 837 q1672 q1673
XSPLIT838 LSmitll_SPLIT 838 q1674 q1675
XSPLIT839 LSmitll_SPLIT 839 q1676 q1677
XSPLIT840 LSmitll_SPLIT 840 q1678 q1679
XSPLIT841 LSmitll_SPLIT 841 q1680 q1681
XSPLIT842 LSmitll_SPLIT 842 q1682 q1683
XSPLIT843 LSmitll_SPLIT 843 q1684 q1685
XSPLIT844 LSmitll_SPLIT 844 q1686 q1687
XSPLIT845 LSmitll_SPLIT 845 q1688 q1689
XSPLIT846 LSmitll_SPLIT 846 q1690 q1691
XSPLIT847 LSmitll_SPLIT 847 q1692 q1693
XSPLIT848 LSmitll_SPLIT 848 q1694 q1695
.ends 1_to_1695_split

