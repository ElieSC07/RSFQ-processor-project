.subckt programmer_instr_memory_final_route program_line4t load4t program_line3t load3t program_line2t load2t program_line1t load1t Addr1_1t Addr1_0t Addr0_1t Addr0_0t read1t read0t read_at_first_addr1t read_at_first_addr0t GCLKt bit_out0 bit_out1 bit_out2 bit_out3 bit_out4 bit_out5 bit_out6

X669 X525-SPLITT-OUT-R-IN X525-SPLITT-OUT-R-INr LSmitll_PTLRX
X670 X525-SPLITT-OUT-R-INr X525-SPLITT-OUT-R-INdc LSmitll_SFQDC
R671 X525-SPLITT-OUT-R-INdc 0 5
X672 X525-SPLITT-OUT-R-IN PAD

X673 X526-SPLITT-OUT-R-IN X526-SPLITT-OUT-R-INr LSmitll_PTLRX
X674 X526-SPLITT-OUT-R-INr X526-SPLITT-OUT-R-INdc LSmitll_SFQDC
R675 X526-SPLITT-OUT-R-INdc 0 5
X676 X526-SPLITT-OUT-R-IN PAD

X677 X527-SPLITT-OUT-R-IN X527-SPLITT-OUT-R-INr LSmitll_PTLRX
X678 X527-SPLITT-OUT-R-INr X527-SPLITT-OUT-R-INdc LSmitll_SFQDC
R679 X527-SPLITT-OUT-R-INdc 0 5
X680 X527-SPLITT-OUT-R-IN PAD

X681 X528-SPLITT-OUT-R-IN X528-SPLITT-OUT-R-INr LSmitll_PTLRX
X682 X528-SPLITT-OUT-R-INr X528-SPLITT-OUT-R-INdc LSmitll_SFQDC
R683 X528-SPLITT-OUT-R-INdc 0 5
X684 X528-SPLITT-OUT-R-IN PAD

X685 X529-SPLITT-OUT-R-IN X529-SPLITT-OUT-R-INr LSmitll_PTLRX
X686 X529-SPLITT-OUT-R-INr X529-SPLITT-OUT-R-INdc LSmitll_SFQDC
R687 X529-SPLITT-OUT-R-INdc 0 5
X688 X529-SPLITT-OUT-R-IN PAD

X689 X530-SPLITT-OUT-R-IN X530-SPLITT-OUT-R-INr LSmitll_PTLRX
X690 X530-SPLITT-OUT-R-INr X530-SPLITT-OUT-R-INdc LSmitll_SFQDC
R691 X530-SPLITT-OUT-R-INdc 0 5
X692 X530-SPLITT-OUT-R-IN PAD

X693 X531-SPLITT-OUT-R-IN X531-SPLITT-OUT-R-INr LSmitll_PTLRX
X694 X531-SPLITT-OUT-R-INr X531-SPLITT-OUT-R-INdc LSmitll_SFQDC
R695 X531-SPLITT-OUT-R-INdc 0 5
X696 X531-SPLITT-OUT-R-IN PAD

X697 X532-SPLITT-OUT-R-IN X532-SPLITT-OUT-R-INr LSmitll_PTLRX
X698 X532-SPLITT-OUT-R-INr X532-SPLITT-OUT-R-INdc LSmitll_SFQDC
R699 X532-SPLITT-OUT-R-INdc 0 5
X700 X532-SPLITT-OUT-R-IN PAD

X701 X533-SPLITT-OUT-R-IN X533-SPLITT-OUT-R-INr LSmitll_PTLRX
X702 X533-SPLITT-OUT-R-INr X533-SPLITT-OUT-R-INdc LSmitll_SFQDC
R703 X533-SPLITT-OUT-R-INdc 0 5
X704 X533-SPLITT-OUT-R-IN PAD

X705 X534-SPLITT-OUT-R-IN X534-SPLITT-OUT-R-INr LSmitll_PTLRX
X706 X534-SPLITT-OUT-R-INr X534-SPLITT-OUT-R-INdc LSmitll_SFQDC
R707 X534-SPLITT-OUT-R-INdc 0 5
X708 X534-SPLITT-OUT-R-IN PAD

X709 X535-SPLITT-OUT-R-IN X535-SPLITT-OUT-R-INr LSmitll_PTLRX
X710 X535-SPLITT-OUT-R-INr X535-SPLITT-OUT-R-INdc LSmitll_SFQDC
R711 X535-SPLITT-OUT-R-INdc 0 5
X712 X535-SPLITT-OUT-R-IN PAD

X713 X536-SPLITT-OUT-R-IN X536-SPLITT-OUT-R-INr LSmitll_PTLRX
X714 X536-SPLITT-OUT-R-INr X536-SPLITT-OUT-R-INdc LSmitll_SFQDC
R715 X536-SPLITT-OUT-R-INdc 0 5
X716 X536-SPLITT-OUT-R-IN PAD

X717 X537-SPLITT-OUT-R-IN X537-SPLITT-OUT-R-INr LSmitll_PTLRX
X718 X537-SPLITT-OUT-R-INr X537-SPLITT-OUT-R-INdc LSmitll_SFQDC
R719 X537-SPLITT-OUT-R-INdc 0 5
X720 X537-SPLITT-OUT-R-IN PAD

X721 X538-SPLITT-OUT-R-IN X538-SPLITT-OUT-R-INr LSmitll_PTLRX
X722 X538-SPLITT-OUT-R-INr X538-SPLITT-OUT-R-INdc LSmitll_SFQDC
R723 X538-SPLITT-OUT-R-INdc 0 5
X724 X538-SPLITT-OUT-R-IN PAD

X725 X539-SPLITT-OUT-R-IN X539-SPLITT-OUT-R-INr LSmitll_PTLRX
X726 X539-SPLITT-OUT-R-INr X539-SPLITT-OUT-R-INdc LSmitll_SFQDC
R727 X539-SPLITT-OUT-R-INdc 0 5
X728 X539-SPLITT-OUT-R-IN PAD

X729 X540-SPLITT-OUT-R-IN X540-SPLITT-OUT-R-INr LSmitll_PTLRX
X730 X540-SPLITT-OUT-R-INr X540-SPLITT-OUT-R-INdc LSmitll_SFQDC
R731 X540-SPLITT-OUT-R-INdc 0 5
X732 X540-SPLITT-OUT-R-IN PAD

X733 X541-SPLITT-OUT-R-IN X541-SPLITT-OUT-R-INr LSmitll_PTLRX
X734 X541-SPLITT-OUT-R-INr X541-SPLITT-OUT-R-INdc LSmitll_SFQDC
R735 X541-SPLITT-OUT-R-INdc 0 5
X736 X541-SPLITT-OUT-R-IN PAD

X737 X542-SPLITT-OUT-R-IN X542-SPLITT-OUT-R-INr LSmitll_PTLRX
X738 X542-SPLITT-OUT-R-INr X542-SPLITT-OUT-R-INdc LSmitll_SFQDC
R739 X542-SPLITT-OUT-R-INdc 0 5
X740 X542-SPLITT-OUT-R-IN PAD

X741 X543-SPLITT-OUT-R-IN X543-SPLITT-OUT-R-INr LSmitll_PTLRX
X742 X543-SPLITT-OUT-R-INr X543-SPLITT-OUT-R-INdc LSmitll_SFQDC
R743 X543-SPLITT-OUT-R-INdc 0 5
X744 X543-SPLITT-OUT-R-IN PAD

X745 X544-SPLITT-OUT-R-IN X544-SPLITT-OUT-R-INr LSmitll_PTLRX
X746 X544-SPLITT-OUT-R-INr X544-SPLITT-OUT-R-INdc LSmitll_SFQDC
R747 X544-SPLITT-OUT-R-INdc 0 5
X748 X544-SPLITT-OUT-R-IN PAD

X749 X545-SPLITT-OUT-R-IN X545-SPLITT-OUT-R-INr LSmitll_PTLRX
X750 X545-SPLITT-OUT-R-INr X545-SPLITT-OUT-R-INdc LSmitll_SFQDC
R751 X545-SPLITT-OUT-R-INdc 0 5
X752 X545-SPLITT-OUT-R-IN PAD

X753 X546-SPLITT-OUT-R-IN X546-SPLITT-OUT-R-INr LSmitll_PTLRX
X754 X546-SPLITT-OUT-R-INr X546-SPLITT-OUT-R-INdc LSmitll_SFQDC
R755 X546-SPLITT-OUT-R-INdc 0 5
X756 X546-SPLITT-OUT-R-IN PAD

X757 X547-SPLITT-OUT-R-IN X547-SPLITT-OUT-R-INr LSmitll_PTLRX
X758 X547-SPLITT-OUT-R-INr X547-SPLITT-OUT-R-INdc LSmitll_SFQDC
R759 X547-SPLITT-OUT-R-INdc 0 5
X760 X547-SPLITT-OUT-R-IN PAD

X761 X548-SPLITT-OUT-R-IN X548-SPLITT-OUT-R-INr LSmitll_PTLRX
X762 X548-SPLITT-OUT-R-INr X548-SPLITT-OUT-R-INdc LSmitll_SFQDC
R763 X548-SPLITT-OUT-R-INdc 0 5
X764 X548-SPLITT-OUT-R-IN PAD

X765 X549-SPLITT-OUT-R-IN X549-SPLITT-OUT-R-INr LSmitll_PTLRX
X766 X549-SPLITT-OUT-R-INr X549-SPLITT-OUT-R-INdc LSmitll_SFQDC
R767 X549-SPLITT-OUT-R-INdc 0 5
X768 X549-SPLITT-OUT-R-IN PAD

X769 X550-SPLITT-OUT-R-IN X550-SPLITT-OUT-R-INr LSmitll_PTLRX
X770 X550-SPLITT-OUT-R-INr X550-SPLITT-OUT-R-INdc LSmitll_SFQDC
R771 X550-SPLITT-OUT-R-INdc 0 5
X772 X550-SPLITT-OUT-R-IN PAD

X773 X551-SPLITT-OUT-R-IN X551-SPLITT-OUT-R-INr LSmitll_PTLRX
X774 X551-SPLITT-OUT-R-INr X551-SPLITT-OUT-R-INdc LSmitll_SFQDC
R775 X551-SPLITT-OUT-R-INdc 0 5
X776 X551-SPLITT-OUT-R-IN PAD

X777 X552-SPLITT-OUT-R-IN X552-SPLITT-OUT-R-INr LSmitll_PTLRX
X778 X552-SPLITT-OUT-R-INr X552-SPLITT-OUT-R-INdc LSmitll_SFQDC
R779 X552-SPLITT-OUT-R-INdc 0 5
X780 X552-SPLITT-OUT-R-IN PAD

X781 X553-SPLITT-OUT-R-IN X553-SPLITT-OUT-R-INr LSmitll_PTLRX
X782 X553-SPLITT-OUT-R-INr X553-SPLITT-OUT-R-INdc LSmitll_SFQDC
R783 X553-SPLITT-OUT-R-INdc 0 5
X784 X553-SPLITT-OUT-R-IN PAD

X785 X554-SPLITT-OUT-R-IN X554-SPLITT-OUT-R-INr LSmitll_PTLRX
X786 X554-SPLITT-OUT-R-INr X554-SPLITT-OUT-R-INdc LSmitll_SFQDC
R787 X554-SPLITT-OUT-R-INdc 0 5
X788 X554-SPLITT-OUT-R-IN PAD

X789 X555-SPLITT-OUT-R-IN X555-SPLITT-OUT-R-INr LSmitll_PTLRX
X790 X555-SPLITT-OUT-R-INr X555-SPLITT-OUT-R-INdc LSmitll_SFQDC
R791 X555-SPLITT-OUT-R-INdc 0 5
X792 X555-SPLITT-OUT-R-IN PAD

X793 X556-SPLITT-OUT-R-IN X556-SPLITT-OUT-R-INr LSmitll_PTLRX
X794 X556-SPLITT-OUT-R-INr X556-SPLITT-OUT-R-INdc LSmitll_SFQDC
R795 X556-SPLITT-OUT-R-INdc 0 5
X796 X556-SPLITT-OUT-R-IN PAD

X797 X557-SPLITT-OUT-R-IN X557-SPLITT-OUT-R-INr LSmitll_PTLRX
X798 X557-SPLITT-OUT-R-INr X557-SPLITT-OUT-R-INdc LSmitll_SFQDC
R799 X557-SPLITT-OUT-R-INdc 0 5
X800 X557-SPLITT-OUT-R-IN PAD

X801 X558-SPLITT-OUT-R-IN X558-SPLITT-OUT-R-INr LSmitll_PTLRX
X802 X558-SPLITT-OUT-R-INr X558-SPLITT-OUT-R-INdc LSmitll_SFQDC
R803 X558-SPLITT-OUT-R-INdc 0 5
X804 X558-SPLITT-OUT-R-IN PAD

X805 X559-SPLITT-OUT-R-IN X559-SPLITT-OUT-R-INr LSmitll_PTLRX
X806 X559-SPLITT-OUT-R-INr X559-SPLITT-OUT-R-INdc LSmitll_SFQDC
R807 X559-SPLITT-OUT-R-INdc 0 5
X808 X559-SPLITT-OUT-R-IN PAD

X809 X560-SPLITT-OUT-R-IN X560-SPLITT-OUT-R-INr LSmitll_PTLRX
X810 X560-SPLITT-OUT-R-INr X560-SPLITT-OUT-R-INdc LSmitll_SFQDC
R811 X560-SPLITT-OUT-R-INdc 0 5
X812 X560-SPLITT-OUT-R-IN PAD

X813 X561-SPLITT-OUT-R-IN X561-SPLITT-OUT-R-INr LSmitll_PTLRX
X814 X561-SPLITT-OUT-R-INr X561-SPLITT-OUT-R-INdc LSmitll_SFQDC
R815 X561-SPLITT-OUT-R-INdc 0 5
X816 X561-SPLITT-OUT-R-IN PAD

X817 X562-SPLITT-OUT-R-IN X562-SPLITT-OUT-R-INr LSmitll_PTLRX
X818 X562-SPLITT-OUT-R-INr X562-SPLITT-OUT-R-INdc LSmitll_SFQDC
R819 X562-SPLITT-OUT-R-INdc 0 5
X820 X562-SPLITT-OUT-R-IN PAD

X821 X563-SPLITT-OUT-R-IN X563-SPLITT-OUT-R-INr LSmitll_PTLRX
X822 X563-SPLITT-OUT-R-INr X563-SPLITT-OUT-R-INdc LSmitll_SFQDC
R823 X563-SPLITT-OUT-R-INdc 0 5
X824 X563-SPLITT-OUT-R-IN PAD

X825 X564-SPLITT-OUT-R-IN X564-SPLITT-OUT-R-INr LSmitll_PTLRX
X826 X564-SPLITT-OUT-R-INr X564-SPLITT-OUT-R-INdc LSmitll_SFQDC
R827 X564-SPLITT-OUT-R-INdc 0 5
X828 X564-SPLITT-OUT-R-IN PAD

X829 X565-SPLITT-OUT-R-IN X565-SPLITT-OUT-R-INr LSmitll_PTLRX
X830 X565-SPLITT-OUT-R-INr X565-SPLITT-OUT-R-INdc LSmitll_SFQDC
R831 X565-SPLITT-OUT-R-INdc 0 5
X832 X565-SPLITT-OUT-R-IN PAD

X833 X566-SPLITT-OUT-R-IN X566-SPLITT-OUT-R-INr LSmitll_PTLRX
X834 X566-SPLITT-OUT-R-INr X566-SPLITT-OUT-R-INdc LSmitll_SFQDC
R835 X566-SPLITT-OUT-R-INdc 0 5
X836 X566-SPLITT-OUT-R-IN PAD

X837 X567-SPLITT-OUT-R-IN X567-SPLITT-OUT-R-INr LSmitll_PTLRX
X838 X567-SPLITT-OUT-R-INr X567-SPLITT-OUT-R-INdc LSmitll_SFQDC
R839 X567-SPLITT-OUT-R-INdc 0 5
X840 X567-SPLITT-OUT-R-IN PAD

X841 X568-SPLITT-OUT-R-IN X568-SPLITT-OUT-R-INr LSmitll_PTLRX
X842 X568-SPLITT-OUT-R-INr X568-SPLITT-OUT-R-INdc LSmitll_SFQDC
R843 X568-SPLITT-OUT-R-INdc 0 5
X844 X568-SPLITT-OUT-R-IN PAD

X845 X569-SPLITT-OUT-R-IN X569-SPLITT-OUT-R-INr LSmitll_PTLRX
X846 X569-SPLITT-OUT-R-INr X569-SPLITT-OUT-R-INdc LSmitll_SFQDC
R847 X569-SPLITT-OUT-R-INdc 0 5
X848 X569-SPLITT-OUT-R-IN PAD

X849 X570-SPLITT-OUT-R-IN X570-SPLITT-OUT-R-INr LSmitll_PTLRX
X850 X570-SPLITT-OUT-R-INr X570-SPLITT-OUT-R-INdc LSmitll_SFQDC
R851 X570-SPLITT-OUT-R-INdc 0 5
X852 X570-SPLITT-OUT-R-IN PAD

X853 X571-SPLITT-OUT-R-IN X571-SPLITT-OUT-R-INr LSmitll_PTLRX
X854 X571-SPLITT-OUT-R-INr X571-SPLITT-OUT-R-INdc LSmitll_SFQDC
R855 X571-SPLITT-OUT-R-INdc 0 5
X856 X571-SPLITT-OUT-R-IN PAD

X857 X572-SPLITT-OUT-R-IN X572-SPLITT-OUT-R-INr LSmitll_PTLRX
X858 X572-SPLITT-OUT-R-INr X572-SPLITT-OUT-R-INdc LSmitll_SFQDC
R859 X572-SPLITT-OUT-R-INdc 0 5
X860 X572-SPLITT-OUT-R-IN PAD

X861 X573-SPLITT-OUT-R-IN X573-SPLITT-OUT-R-INr LSmitll_PTLRX
X862 X573-SPLITT-OUT-R-INr X573-SPLITT-OUT-R-INdc LSmitll_SFQDC
R863 X573-SPLITT-OUT-R-INdc 0 5
X864 X573-SPLITT-OUT-R-IN PAD

X865 X574-SPLITT-OUT-R-IN X574-SPLITT-OUT-R-INr LSmitll_PTLRX
X866 X574-SPLITT-OUT-R-INr X574-SPLITT-OUT-R-INdc LSmitll_SFQDC
R867 X574-SPLITT-OUT-R-INdc 0 5
X868 X574-SPLITT-OUT-R-IN PAD

X869 X575-SPLITT-OUT-R-IN X575-SPLITT-OUT-R-INr LSmitll_PTLRX
X870 X575-SPLITT-OUT-R-INr X575-SPLITT-OUT-R-INdc LSmitll_SFQDC
R871 X575-SPLITT-OUT-R-INdc 0 5
X872 X575-SPLITT-OUT-R-IN PAD

t877 X1-LSmitll_SPLITT-OUT-X189-LSmitll_SPLITT-INt 0 X1-LSmitll_SPLITT-OUT-X189-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t878 X1-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-INt 0 X1-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-IN 0 z0=5 td=4.1ps
X1 load1 X1-LSmitll_SPLITT-OUT-X189-LSmitll_SPLITT-INt X1-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-INt LSmitll_SPLITT

t879 X2-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-INt 0 X2-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t880 X2-LSmitll_SPLITT-OUT-X17-LSmitll_DFFT-INt 0 X2-LSmitll_SPLITT-OUT-X17-LSmitll_DFFT-IN 0 z0=5 td=4.1ps
X2 program_line1 X2-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-INt X2-LSmitll_SPLITT-OUT-X17-LSmitll_DFFT-INt LSmitll_SPLITT

t881 X3-LSmitll_SPLITT-OUT-X196-LSmitll_SPLITT-INt 0 X3-LSmitll_SPLITT-OUT-X196-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t882 X3-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-INt 0 X3-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-IN 0 z0=5 td=4.0ps
X3 load2 X3-LSmitll_SPLITT-OUT-X196-LSmitll_SPLITT-INt X3-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-INt LSmitll_SPLITT

t883 X4-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-INt 0 X4-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t884 X4-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-INt 0 X4-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-IN 0 z0=5 td=5.2ps
X4 program_line2 X4-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-INt X4-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-INt LSmitll_SPLITT

t885 X5-LSmitll_SPLITT-OUT-X203-LSmitll_SPLITT-INt 0 X5-LSmitll_SPLITT-OUT-X203-LSmitll_SPLITT-IN 0 z0=5 td=4.6ps
t886 X5-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-INt 0 X5-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X5 load3 X5-LSmitll_SPLITT-OUT-X203-LSmitll_SPLITT-INt X5-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-INt LSmitll_SPLITT

t887 X6-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-INt 0 X6-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t888 X6-LSmitll_SPLITT-OUT-X23-LSmitll_DFFT-INt 0 X6-LSmitll_SPLITT-OUT-X23-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X6 program_line3 X6-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-INt X6-LSmitll_SPLITT-OUT-X23-LSmitll_DFFT-INt LSmitll_SPLITT

t889 X7-LSmitll_SPLITT-OUT-X210-LSmitll_SPLITT-INt 0 X7-LSmitll_SPLITT-OUT-X210-LSmitll_SPLITT-IN 0 z0=5 td=9.8ps
t890 X7-LSmitll_SPLITT-OUT-X27-LSmitll_DFFT-INt 0 X7-LSmitll_SPLITT-OUT-X27-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X7 load4 X7-LSmitll_SPLITT-OUT-X210-LSmitll_SPLITT-INt X7-LSmitll_SPLITT-OUT-X27-LSmitll_DFFT-INt LSmitll_SPLITT

t891 X8-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-INt 0 X8-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-IN 0 z0=5 td=2.6ps
t892 X8-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-INt 0 X8-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X8 program_line4 X8-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-INt X8-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-INt LSmitll_SPLITT

t893 X9-LSmitll_SPLITT-OUT-X37-LSmitll_NOTT-INt 0 X9-LSmitll_SPLITT-OUT-X37-LSmitll_NOTT-IN 0 z0=5 td=1.2ps
t894 X9-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-INt 0 X9-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X9 Addr1_0 X9-LSmitll_SPLITT-OUT-X37-LSmitll_NOTT-INt X9-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-INt LSmitll_SPLITT

t895 X10-LSmitll_SPLITT-OUT-X38-LSmitll_NOTT-INt 0 X10-LSmitll_SPLITT-OUT-X38-LSmitll_NOTT-IN 0 z0=5 td=4.7ps
t896 X10-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-INt 0 X10-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-IN 0 z0=5 td=6.3ps
X10 Addr0_0 X10-LSmitll_SPLITT-OUT-X38-LSmitll_NOTT-INt X10-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-INt LSmitll_SPLITT

t897 X11-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-INt 0 X11-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-IN 0 z0=5 td=1.2ps
t898 X11-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-INt 0 X11-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-IN 0 z0=5 td=4.9ps
X11 read_at_first_addr0 X11-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-INt X11-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-INt LSmitll_SPLITT

t899 X12-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-INt 0 X12-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-IN 0 z0=5 td=4.0ps
t900 X12-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-INt 0 X12-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-IN 0 z0=5 td=2.1ps
X12 read0 X12-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-INt X12-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-INt LSmitll_SPLITT

t901 X13-LSmitll_SPLITT-OUT-X39-LSmitll_NOTT-INt 0 X13-LSmitll_SPLITT-OUT-X39-LSmitll_NOTT-IN 0 z0=5 td=5.9ps
t902 X13-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-INt 0 X13-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-IN 0 z0=5 td=4.9ps
X13 Addr1_1 X13-LSmitll_SPLITT-OUT-X39-LSmitll_NOTT-INt X13-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-INt LSmitll_SPLITT

t903 X14-LSmitll_SPLITT-OUT-X40-LSmitll_NOTT-INt 0 X14-LSmitll_SPLITT-OUT-X40-LSmitll_NOTT-IN 0 z0=5 td=1.2ps
t904 X14-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-INt 0 X14-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
X14 Addr0_1 X14-LSmitll_SPLITT-OUT-X40-LSmitll_NOTT-INt X14-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-INt LSmitll_SPLITT

t905 X15-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-INt 0 X15-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-IN 0 z0=5 td=1.7ps
t906 X15-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-INt 0 X15-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-IN 0 z0=5 td=1.4ps
X15 read_at_first_addr1 X15-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-INt X15-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-INt LSmitll_SPLITT

t907 X16-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-INt 0 X16-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-IN 0 z0=5 td=1.8ps
t908 X16-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-INt 0 X16-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-IN 0 z0=5 td=2.3ps
X16 read1 X16-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-INt X16-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-INt LSmitll_SPLITT

t909 X17-LSmitll_DFFT-OUT-X41-LSmitll_SPLITT-INt 0 X17-LSmitll_DFFT-OUT-X41-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
X17 X2-LSmitll_SPLITT-OUT-X17-LSmitll_DFFT-IN X450-LSmitll_SPLITT-OUT-X17-LSmitll_DFFT-IN X17-LSmitll_DFFT-OUT-X41-LSmitll_SPLITT-INt LSmitll_DFFT

t910 X18-LSmitll_DFFT-OUT-X19-LSmitll_DFFT-INt 0 X18-LSmitll_DFFT-OUT-X19-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X18 X1-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-IN X455-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-IN X18-LSmitll_DFFT-OUT-X19-LSmitll_DFFT-INt LSmitll_DFFT

t911 X19-LSmitll_DFFT-OUT-X42-LSmitll_SPLITT-INt 0 X19-LSmitll_DFFT-OUT-X42-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X19 X18-LSmitll_DFFT-OUT-X19-LSmitll_DFFT-IN X525-LSmitll_SPLITT-OUT-X19-LSmitll_DFFT-IN X19-LSmitll_DFFT-OUT-X42-LSmitll_SPLITT-INt LSmitll_DFFT

t912 X20-LSmitll_DFFT-OUT-X43-LSmitll_SPLITT-INt 0 X20-LSmitll_DFFT-OUT-X43-LSmitll_SPLITT-IN 0 z0=5 td=6.5ps
X20 X4-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-IN X425-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-IN X20-LSmitll_DFFT-OUT-X43-LSmitll_SPLITT-INt LSmitll_DFFT

t913 X21-LSmitll_DFFT-OUT-X22-LSmitll_DFFT-INt 0 X21-LSmitll_DFFT-OUT-X22-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X21 X3-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-IN X432-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-IN X21-LSmitll_DFFT-OUT-X22-LSmitll_DFFT-INt LSmitll_DFFT

t914 X22-LSmitll_DFFT-OUT-X44-LSmitll_SPLITT-INt 0 X22-LSmitll_DFFT-OUT-X44-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
X22 X21-LSmitll_DFFT-OUT-X22-LSmitll_DFFT-IN X430-LSmitll_SPLITT-OUT-X22-LSmitll_DFFT-IN X22-LSmitll_DFFT-OUT-X44-LSmitll_SPLITT-INt LSmitll_DFFT

t915 X23-LSmitll_DFFT-OUT-X45-LSmitll_SPLITT-INt 0 X23-LSmitll_DFFT-OUT-X45-LSmitll_SPLITT-IN 0 z0=5 td=18.7ps
X23 X6-LSmitll_SPLITT-OUT-X23-LSmitll_DFFT-IN X430-LSmitll_SPLITT-OUT-X23-LSmitll_DFFT-IN X23-LSmitll_DFFT-OUT-X45-LSmitll_SPLITT-INt LSmitll_DFFT

t916 X24-LSmitll_DFFT-OUT-X25-LSmitll_DFFT-INt 0 X24-LSmitll_DFFT-OUT-X25-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X24 X5-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-IN X348-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-IN X24-LSmitll_DFFT-OUT-X25-LSmitll_DFFT-INt LSmitll_DFFT

t917 X25-LSmitll_DFFT-OUT-X46-LSmitll_SPLITT-INt 0 X25-LSmitll_DFFT-OUT-X46-LSmitll_SPLITT-IN 0 z0=5 td=11.2ps
X25 X24-LSmitll_DFFT-OUT-X25-LSmitll_DFFT-IN X353-LSmitll_SPLITT-OUT-X25-LSmitll_DFFT-IN X25-LSmitll_DFFT-OUT-X46-LSmitll_SPLITT-INt LSmitll_DFFT

t918 X26-LSmitll_DFFT-OUT-X47-LSmitll_SPLITT-INt 0 X26-LSmitll_DFFT-OUT-X47-LSmitll_SPLITT-IN 0 z0=5 td=5.7ps
X26 X8-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-IN X323-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-IN X26-LSmitll_DFFT-OUT-X47-LSmitll_SPLITT-INt LSmitll_DFFT

t919 X27-LSmitll_DFFT-OUT-X28-LSmitll_DFFT-INt 0 X27-LSmitll_DFFT-OUT-X28-LSmitll_DFFT-IN 0 z0=5 td=4.5ps
X27 X7-LSmitll_SPLITT-OUT-X27-LSmitll_DFFT-IN X328-LSmitll_SPLITT-OUT-X27-LSmitll_DFFT-IN X27-LSmitll_DFFT-OUT-X28-LSmitll_DFFT-INt LSmitll_DFFT

t920 X28-LSmitll_DFFT-OUT-X48-LSmitll_SPLITT-INt 0 X28-LSmitll_DFFT-OUT-X48-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X28 X27-LSmitll_DFFT-OUT-X28-LSmitll_DFFT-IN X323-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-IN X28-LSmitll_DFFT-OUT-X48-LSmitll_SPLITT-INt LSmitll_DFFT

t921 X29-LSmitll_DFFT-OUT-X65-LSmitll_AND2T-INt 0 X29-LSmitll_DFFT-OUT-X65-LSmitll_AND2T-IN 0 z0=5 td=9.7ps
X29 X9-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-IN X442-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-IN X29-LSmitll_DFFT-OUT-X65-LSmitll_AND2T-INt LSmitll_DFFT

t922 X30-LSmitll_DFFT-OUT-X67-LSmitll_AND2T-INt 0 X30-LSmitll_DFFT-OUT-X67-LSmitll_AND2T-IN 0 z0=5 td=3.6ps
X30 X10-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-IN X374-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-IN X30-LSmitll_DFFT-OUT-X67-LSmitll_AND2T-INt LSmitll_DFFT

t923 X31-LSmitll_DFFT-OUT-X69-LSmitll_AND2T-INt 0 X31-LSmitll_DFFT-OUT-X69-LSmitll_AND2T-IN 0 z0=5 td=5.6ps
X31 X13-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-IN X388-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-IN X31-LSmitll_DFFT-OUT-X69-LSmitll_AND2T-INt LSmitll_DFFT

t924 X32-LSmitll_DFFT-OUT-X71-LSmitll_AND2T-INt 0 X32-LSmitll_DFFT-OUT-X71-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X32 X14-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-IN X518-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-IN X32-LSmitll_DFFT-OUT-X71-LSmitll_AND2T-INt LSmitll_DFFT

t925 X33-LSmitll_OR2T-OUT-X49-LSmitll_SPLITT-INt 0 X33-LSmitll_OR2T-OUT-X49-LSmitll_SPLITT-IN 0 z0=5 td=16.3ps
X33 X11-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-IN X12-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-IN X526-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-IN X33-LSmitll_OR2T-OUT-X49-LSmitll_SPLITT-INt LSmitll_OR2T

t926 X34-LSmitll_OR2T-OUT-X50-LSmitll_SPLITT-INt 0 X34-LSmitll_OR2T-OUT-X50-LSmitll_SPLITT-IN 0 z0=5 td=12.3ps
X34 X11-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-IN X12-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-IN X412-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-IN X34-LSmitll_OR2T-OUT-X50-LSmitll_SPLITT-INt LSmitll_OR2T

t927 X35-LSmitll_OR2T-OUT-X51-LSmitll_SPLITT-INt 0 X35-LSmitll_OR2T-OUT-X51-LSmitll_SPLITT-IN 0 z0=5 td=12.6ps
X35 X15-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-IN X16-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-IN X489-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-IN X35-LSmitll_OR2T-OUT-X51-LSmitll_SPLITT-INt LSmitll_OR2T

t928 X36-LSmitll_OR2T-OUT-X52-LSmitll_SPLITT-INt 0 X36-LSmitll_OR2T-OUT-X52-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
X36 X15-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-IN X16-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-IN X494-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-IN X36-LSmitll_OR2T-OUT-X52-LSmitll_SPLITT-INt LSmitll_OR2T

t929 X37-LSmitll_NOTT-OUT-X66-LSmitll_AND2T-INt 0 X37-LSmitll_NOTT-OUT-X66-LSmitll_AND2T-IN 0 z0=5 td=4.6ps
X37 X9-LSmitll_SPLITT-OUT-X37-LSmitll_NOTT-IN X427-LSmitll_SPLITT-OUT-X37-LSmitll_NOTT-IN X37-LSmitll_NOTT-OUT-X66-LSmitll_AND2T-INt LSmitll_NOTT

t930 X38-LSmitll_NOTT-OUT-X68-LSmitll_AND2T-INt 0 X38-LSmitll_NOTT-OUT-X68-LSmitll_AND2T-IN 0 z0=5 td=5.5ps
X38 X10-LSmitll_SPLITT-OUT-X38-LSmitll_NOTT-IN X527-LSmitll_SPLITT-OUT-X38-LSmitll_NOTT-IN X38-LSmitll_NOTT-OUT-X68-LSmitll_AND2T-INt LSmitll_NOTT

t931 X39-LSmitll_NOTT-OUT-X70-LSmitll_AND2T-INt 0 X39-LSmitll_NOTT-OUT-X70-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
X39 X13-LSmitll_SPLITT-OUT-X39-LSmitll_NOTT-IN X393-LSmitll_SPLITT-OUT-X39-LSmitll_NOTT-IN X39-LSmitll_NOTT-OUT-X70-LSmitll_AND2T-INt LSmitll_NOTT

t932 X40-LSmitll_NOTT-OUT-X72-LSmitll_AND2T-INt 0 X40-LSmitll_NOTT-OUT-X72-LSmitll_AND2T-IN 0 z0=5 td=4.3ps
X40 X14-LSmitll_SPLITT-OUT-X40-LSmitll_NOTT-IN X528-LSmitll_SPLITT-OUT-X40-LSmitll_NOTT-IN X40-LSmitll_NOTT-OUT-X72-LSmitll_AND2T-INt LSmitll_NOTT

t933 X41-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-INt 0 X41-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t934 X41-LSmitll_SPLITT-OUT-X53-LSmitll_DFFT-INt 0 X41-LSmitll_SPLITT-OUT-X53-LSmitll_DFFT-IN 0 z0=5 td=3.0ps
X41 X17-LSmitll_DFFT-OUT-X41-LSmitll_SPLITT-IN X41-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-INt X41-LSmitll_SPLITT-OUT-X53-LSmitll_DFFT-INt LSmitll_SPLITT

t935 X42-LSmitll_SPLITT-OUT-X190-LSmitll_SPLITT-INt 0 X42-LSmitll_SPLITT-OUT-X190-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t936 X42-LSmitll_SPLITT-OUT-X54-LSmitll_DFFT-INt 0 X42-LSmitll_SPLITT-OUT-X54-LSmitll_DFFT-IN 0 z0=5 td=2.7ps
X42 X19-LSmitll_DFFT-OUT-X42-LSmitll_SPLITT-IN X42-LSmitll_SPLITT-OUT-X190-LSmitll_SPLITT-INt X42-LSmitll_SPLITT-OUT-X54-LSmitll_DFFT-INt LSmitll_SPLITT

t937 X43-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt 0 X43-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t938 X43-LSmitll_SPLITT-OUT-X56-LSmitll_DFFT-INt 0 X43-LSmitll_SPLITT-OUT-X56-LSmitll_DFFT-IN 0 z0=5 td=2.0ps
X43 X20-LSmitll_DFFT-OUT-X43-LSmitll_SPLITT-IN X43-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt X43-LSmitll_SPLITT-OUT-X56-LSmitll_DFFT-INt LSmitll_SPLITT

t939 X44-LSmitll_SPLITT-OUT-X197-LSmitll_SPLITT-INt 0 X44-LSmitll_SPLITT-OUT-X197-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
t940 X44-LSmitll_SPLITT-OUT-X57-LSmitll_DFFT-INt 0 X44-LSmitll_SPLITT-OUT-X57-LSmitll_DFFT-IN 0 z0=5 td=2.9ps
X44 X22-LSmitll_DFFT-OUT-X44-LSmitll_SPLITT-IN X44-LSmitll_SPLITT-OUT-X197-LSmitll_SPLITT-INt X44-LSmitll_SPLITT-OUT-X57-LSmitll_DFFT-INt LSmitll_SPLITT

t941 X45-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-INt 0 X45-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-IN 0 z0=5 td=3.9ps
t942 X45-LSmitll_SPLITT-OUT-X59-LSmitll_DFFT-INt 0 X45-LSmitll_SPLITT-OUT-X59-LSmitll_DFFT-IN 0 z0=5 td=2.7ps
X45 X23-LSmitll_DFFT-OUT-X45-LSmitll_SPLITT-IN X45-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-INt X45-LSmitll_SPLITT-OUT-X59-LSmitll_DFFT-INt LSmitll_SPLITT

t943 X46-LSmitll_SPLITT-OUT-X204-LSmitll_SPLITT-INt 0 X46-LSmitll_SPLITT-OUT-X204-LSmitll_SPLITT-IN 0 z0=5 td=4.8ps
t944 X46-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-INt 0 X46-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-IN 0 z0=5 td=2.5ps
X46 X25-LSmitll_DFFT-OUT-X46-LSmitll_SPLITT-IN X46-LSmitll_SPLITT-OUT-X204-LSmitll_SPLITT-INt X46-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-INt LSmitll_SPLITT

t945 X47-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-INt 0 X47-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t946 X47-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-INt 0 X47-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-IN 0 z0=5 td=4.9ps
X47 X26-LSmitll_DFFT-OUT-X47-LSmitll_SPLITT-IN X47-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-INt X47-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-INt LSmitll_SPLITT

t947 X48-LSmitll_SPLITT-OUT-X211-LSmitll_SPLITT-INt 0 X48-LSmitll_SPLITT-OUT-X211-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
t948 X48-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-INt 0 X48-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-IN 0 z0=5 td=2.8ps
X48 X28-LSmitll_DFFT-OUT-X48-LSmitll_SPLITT-IN X48-LSmitll_SPLITT-OUT-X211-LSmitll_SPLITT-INt X48-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-INt LSmitll_SPLITT

t949 X49-LSmitll_SPLITT-OUT-X66-LSmitll_AND2T-INt 0 X49-LSmitll_SPLITT-OUT-X66-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
t950 X49-LSmitll_SPLITT-OUT-X65-LSmitll_AND2T-INt 0 X49-LSmitll_SPLITT-OUT-X65-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X49 X33-LSmitll_OR2T-OUT-X49-LSmitll_SPLITT-IN X49-LSmitll_SPLITT-OUT-X66-LSmitll_AND2T-INt X49-LSmitll_SPLITT-OUT-X65-LSmitll_AND2T-INt LSmitll_SPLITT

t951 X50-LSmitll_SPLITT-OUT-X68-LSmitll_AND2T-INt 0 X50-LSmitll_SPLITT-OUT-X68-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t952 X50-LSmitll_SPLITT-OUT-X67-LSmitll_AND2T-INt 0 X50-LSmitll_SPLITT-OUT-X67-LSmitll_AND2T-IN 0 z0=5 td=2.6ps
X50 X34-LSmitll_OR2T-OUT-X50-LSmitll_SPLITT-IN X50-LSmitll_SPLITT-OUT-X68-LSmitll_AND2T-INt X50-LSmitll_SPLITT-OUT-X67-LSmitll_AND2T-INt LSmitll_SPLITT

t953 X51-LSmitll_SPLITT-OUT-X70-LSmitll_AND2T-INt 0 X51-LSmitll_SPLITT-OUT-X70-LSmitll_AND2T-IN 0 z0=5 td=4.9ps
t954 X51-LSmitll_SPLITT-OUT-X69-LSmitll_AND2T-INt 0 X51-LSmitll_SPLITT-OUT-X69-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X51 X35-LSmitll_OR2T-OUT-X51-LSmitll_SPLITT-IN X51-LSmitll_SPLITT-OUT-X70-LSmitll_AND2T-INt X51-LSmitll_SPLITT-OUT-X69-LSmitll_AND2T-INt LSmitll_SPLITT

t955 X52-LSmitll_SPLITT-OUT-X72-LSmitll_AND2T-INt 0 X52-LSmitll_SPLITT-OUT-X72-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t956 X52-LSmitll_SPLITT-OUT-X71-LSmitll_AND2T-INt 0 X52-LSmitll_SPLITT-OUT-X71-LSmitll_AND2T-IN 0 z0=5 td=4.1ps
X52 X36-LSmitll_OR2T-OUT-X52-LSmitll_SPLITT-IN X52-LSmitll_SPLITT-OUT-X72-LSmitll_AND2T-INt X52-LSmitll_SPLITT-OUT-X71-LSmitll_AND2T-INt LSmitll_SPLITT

t957 X53-LSmitll_DFFT-OUT-X73-LSmitll_SPLITT-INt 0 X53-LSmitll_DFFT-OUT-X73-LSmitll_SPLITT-IN 0 z0=5 td=3.4ps
X53 X41-LSmitll_SPLITT-OUT-X53-LSmitll_DFFT-IN X457-LSmitll_SPLITT-OUT-X53-LSmitll_DFFT-IN X53-LSmitll_DFFT-OUT-X73-LSmitll_SPLITT-INt LSmitll_DFFT

t958 X54-LSmitll_DFFT-OUT-X55-LSmitll_DFFT-INt 0 X54-LSmitll_DFFT-OUT-X55-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X54 X42-LSmitll_SPLITT-OUT-X54-LSmitll_DFFT-IN X457-LSmitll_SPLITT-OUT-X54-LSmitll_DFFT-IN X54-LSmitll_DFFT-OUT-X55-LSmitll_DFFT-INt LSmitll_DFFT

t959 X55-LSmitll_DFFT-OUT-X74-LSmitll_SPLITT-INt 0 X55-LSmitll_DFFT-OUT-X74-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X55 X54-LSmitll_DFFT-OUT-X55-LSmitll_DFFT-IN X529-LSmitll_SPLITT-OUT-X55-LSmitll_DFFT-IN X55-LSmitll_DFFT-OUT-X74-LSmitll_SPLITT-INt LSmitll_DFFT

t960 X56-LSmitll_DFFT-OUT-X75-LSmitll_SPLITT-INt 0 X56-LSmitll_DFFT-OUT-X75-LSmitll_SPLITT-IN 0 z0=5 td=7.4ps
X56 X43-LSmitll_SPLITT-OUT-X56-LSmitll_DFFT-IN X432-LSmitll_SPLITT-OUT-X56-LSmitll_DFFT-IN X56-LSmitll_DFFT-OUT-X75-LSmitll_SPLITT-INt LSmitll_DFFT

t961 X57-LSmitll_DFFT-OUT-X58-LSmitll_DFFT-INt 0 X57-LSmitll_DFFT-OUT-X58-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X57 X44-LSmitll_SPLITT-OUT-X57-LSmitll_DFFT-IN X452-LSmitll_SPLITT-OUT-X57-LSmitll_DFFT-IN X57-LSmitll_DFFT-OUT-X58-LSmitll_DFFT-INt LSmitll_DFFT

t962 X58-LSmitll_DFFT-OUT-X76-LSmitll_SPLITT-INt 0 X58-LSmitll_DFFT-OUT-X76-LSmitll_SPLITT-IN 0 z0=5 td=4.7ps
X58 X57-LSmitll_DFFT-OUT-X58-LSmitll_DFFT-IN X452-LSmitll_SPLITT-OUT-X58-LSmitll_DFFT-IN X58-LSmitll_DFFT-OUT-X76-LSmitll_SPLITT-INt LSmitll_DFFT

t963 X59-LSmitll_DFFT-OUT-X77-LSmitll_SPLITT-INt 0 X59-LSmitll_DFFT-OUT-X77-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X59 X45-LSmitll_SPLITT-OUT-X59-LSmitll_DFFT-IN X427-LSmitll_SPLITT-OUT-X59-LSmitll_DFFT-IN X59-LSmitll_DFFT-OUT-X77-LSmitll_SPLITT-INt LSmitll_DFFT

t964 X60-LSmitll_DFFT-OUT-X61-LSmitll_DFFT-INt 0 X60-LSmitll_DFFT-OUT-X61-LSmitll_DFFT-IN 0 z0=5 td=2.9ps
X60 X46-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-IN X350-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-IN X60-LSmitll_DFFT-OUT-X61-LSmitll_DFFT-INt LSmitll_DFFT

t965 X61-LSmitll_DFFT-OUT-X78-LSmitll_SPLITT-INt 0 X61-LSmitll_DFFT-OUT-X78-LSmitll_SPLITT-IN 0 z0=5 td=5.1ps
X61 X60-LSmitll_DFFT-OUT-X61-LSmitll_DFFT-IN X359-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-IN X61-LSmitll_DFFT-OUT-X78-LSmitll_SPLITT-INt LSmitll_DFFT

t966 X62-LSmitll_DFFT-OUT-X79-LSmitll_SPLITT-INt 0 X62-LSmitll_DFFT-OUT-X79-LSmitll_SPLITT-IN 0 z0=5 td=9.4ps
X62 X47-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-IN X334-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-IN X62-LSmitll_DFFT-OUT-X79-LSmitll_SPLITT-INt LSmitll_DFFT

t967 X63-LSmitll_DFFT-OUT-X64-LSmitll_DFFT-INt 0 X63-LSmitll_DFFT-OUT-X64-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X63 X48-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-IN X325-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-IN X63-LSmitll_DFFT-OUT-X64-LSmitll_DFFT-INt LSmitll_DFFT

t968 X64-LSmitll_DFFT-OUT-X80-LSmitll_SPLITT-INt 0 X64-LSmitll_DFFT-OUT-X80-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X64 X63-LSmitll_DFFT-OUT-X64-LSmitll_DFFT-IN X325-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-IN X64-LSmitll_DFFT-OUT-X80-LSmitll_SPLITT-INt LSmitll_DFFT

t969 X65-LSmitll_AND2T-OUT-X81-LSmitll_SPLITT-INt 0 X65-LSmitll_AND2T-OUT-X81-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X65 X29-LSmitll_DFFT-OUT-X65-LSmitll_AND2T-IN X49-LSmitll_SPLITT-OUT-X65-LSmitll_AND2T-IN X365-LSmitll_SPLITT-OUT-X65-LSmitll_AND2T-IN X65-LSmitll_AND2T-OUT-X81-LSmitll_SPLITT-INt LSmitll_AND2T

t970 X66-LSmitll_AND2T-OUT-X82-LSmitll_SPLITT-INt 0 X66-LSmitll_AND2T-OUT-X82-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X66 X37-LSmitll_NOTT-OUT-X66-LSmitll_AND2T-IN X49-LSmitll_SPLITT-OUT-X66-LSmitll_AND2T-IN X436-LSmitll_SPLITT-OUT-X66-LSmitll_AND2T-IN X66-LSmitll_AND2T-OUT-X82-LSmitll_SPLITT-INt LSmitll_AND2T

t971 X67-LSmitll_AND2T-OUT-X83-LSmitll_SPLITT-INt 0 X67-LSmitll_AND2T-OUT-X83-LSmitll_SPLITT-IN 0 z0=5 td=9.2ps
X67 X30-LSmitll_DFFT-OUT-X67-LSmitll_AND2T-IN X50-LSmitll_SPLITT-OUT-X67-LSmitll_AND2T-IN X379-LSmitll_SPLITT-OUT-X67-LSmitll_AND2T-IN X67-LSmitll_AND2T-OUT-X83-LSmitll_SPLITT-INt LSmitll_AND2T

t972 X68-LSmitll_AND2T-OUT-X84-LSmitll_SPLITT-INt 0 X68-LSmitll_AND2T-OUT-X84-LSmitll_SPLITT-IN 0 z0=5 td=8.7ps
X68 X38-LSmitll_NOTT-OUT-X68-LSmitll_AND2T-IN X50-LSmitll_SPLITT-OUT-X68-LSmitll_AND2T-IN X530-LSmitll_SPLITT-OUT-X68-LSmitll_AND2T-IN X68-LSmitll_AND2T-OUT-X84-LSmitll_SPLITT-INt LSmitll_AND2T

t973 X69-LSmitll_AND2T-OUT-X85-LSmitll_SPLITT-INt 0 X69-LSmitll_AND2T-OUT-X85-LSmitll_SPLITT-IN 0 z0=5 td=8.8ps
X69 X31-LSmitll_DFFT-OUT-X69-LSmitll_AND2T-IN X51-LSmitll_SPLITT-OUT-X69-LSmitll_AND2T-IN X531-LSmitll_SPLITT-OUT-X69-LSmitll_AND2T-IN X69-LSmitll_AND2T-OUT-X85-LSmitll_SPLITT-INt LSmitll_AND2T

t974 X70-LSmitll_AND2T-OUT-X86-LSmitll_SPLITT-INt 0 X70-LSmitll_AND2T-OUT-X86-LSmitll_SPLITT-IN 0 z0=5 td=8.6ps
X70 X39-LSmitll_NOTT-OUT-X70-LSmitll_AND2T-IN X51-LSmitll_SPLITT-OUT-X70-LSmitll_AND2T-IN X393-LSmitll_SPLITT-OUT-X70-LSmitll_AND2T-IN X70-LSmitll_AND2T-OUT-X86-LSmitll_SPLITT-INt LSmitll_AND2T

t975 X71-LSmitll_AND2T-OUT-X87-LSmitll_SPLITT-INt 0 X71-LSmitll_AND2T-OUT-X87-LSmitll_SPLITT-IN 0 z0=5 td=18.3ps
X71 X32-LSmitll_DFFT-OUT-X71-LSmitll_AND2T-IN X52-LSmitll_SPLITT-OUT-X71-LSmitll_AND2T-IN X532-LSmitll_SPLITT-OUT-X71-LSmitll_AND2T-IN X71-LSmitll_AND2T-OUT-X87-LSmitll_SPLITT-INt LSmitll_AND2T

t976 X72-LSmitll_AND2T-OUT-X88-LSmitll_SPLITT-INt 0 X72-LSmitll_AND2T-OUT-X88-LSmitll_SPLITT-IN 0 z0=5 td=7.8ps
X72 X40-LSmitll_NOTT-OUT-X72-LSmitll_AND2T-IN X52-LSmitll_SPLITT-OUT-X72-LSmitll_AND2T-IN X513-LSmitll_SPLITT-OUT-X72-LSmitll_AND2T-IN X72-LSmitll_AND2T-OUT-X88-LSmitll_SPLITT-INt LSmitll_AND2T

t977 X73-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-INt 0 X73-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
t978 X73-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-INt 0 X73-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-IN 0 z0=5 td=3.4ps
X73 X53-LSmitll_DFFT-OUT-X73-LSmitll_SPLITT-IN X73-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-INt X73-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-INt LSmitll_SPLITT

t979 X74-LSmitll_SPLITT-OUT-X191-LSmitll_SPLITT-INt 0 X74-LSmitll_SPLITT-OUT-X191-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
t980 X74-LSmitll_SPLITT-OUT-X90-LSmitll_DFFT-INt 0 X74-LSmitll_SPLITT-OUT-X90-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
X74 X55-LSmitll_DFFT-OUT-X74-LSmitll_SPLITT-IN X74-LSmitll_SPLITT-OUT-X191-LSmitll_SPLITT-INt X74-LSmitll_SPLITT-OUT-X90-LSmitll_DFFT-INt LSmitll_SPLITT

t981 X75-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-INt 0 X75-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-IN 0 z0=5 td=1.9ps
t982 X75-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-INt 0 X75-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X75 X56-LSmitll_DFFT-OUT-X75-LSmitll_SPLITT-IN X75-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-INt X75-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-INt LSmitll_SPLITT

t983 X76-LSmitll_SPLITT-OUT-X198-LSmitll_SPLITT-INt 0 X76-LSmitll_SPLITT-OUT-X198-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t984 X76-LSmitll_SPLITT-OUT-X93-LSmitll_DFFT-INt 0 X76-LSmitll_SPLITT-OUT-X93-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X76 X58-LSmitll_DFFT-OUT-X76-LSmitll_SPLITT-IN X76-LSmitll_SPLITT-OUT-X198-LSmitll_SPLITT-INt X76-LSmitll_SPLITT-OUT-X93-LSmitll_DFFT-INt LSmitll_SPLITT

t985 X77-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-INt 0 X77-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t986 X77-LSmitll_SPLITT-OUT-X95-LSmitll_DFFT-INt 0 X77-LSmitll_SPLITT-OUT-X95-LSmitll_DFFT-IN 0 z0=5 td=4.6ps
X77 X59-LSmitll_DFFT-OUT-X77-LSmitll_SPLITT-IN X77-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-INt X77-LSmitll_SPLITT-OUT-X95-LSmitll_DFFT-INt LSmitll_SPLITT

t987 X78-LSmitll_SPLITT-OUT-X205-LSmitll_SPLITT-INt 0 X78-LSmitll_SPLITT-OUT-X205-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t988 X78-LSmitll_SPLITT-OUT-X96-LSmitll_DFFT-INt 0 X78-LSmitll_SPLITT-OUT-X96-LSmitll_DFFT-IN 0 z0=5 td=3.9ps
X78 X61-LSmitll_DFFT-OUT-X78-LSmitll_SPLITT-IN X78-LSmitll_SPLITT-OUT-X205-LSmitll_SPLITT-INt X78-LSmitll_SPLITT-OUT-X96-LSmitll_DFFT-INt LSmitll_SPLITT

t989 X79-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-INt 0 X79-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-IN 0 z0=5 td=3.0ps
t990 X79-LSmitll_SPLITT-OUT-X98-LSmitll_DFFT-INt 0 X79-LSmitll_SPLITT-OUT-X98-LSmitll_DFFT-IN 0 z0=5 td=3.0ps
X79 X62-LSmitll_DFFT-OUT-X79-LSmitll_SPLITT-IN X79-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-INt X79-LSmitll_SPLITT-OUT-X98-LSmitll_DFFT-INt LSmitll_SPLITT

t991 X80-LSmitll_SPLITT-OUT-X212-LSmitll_SPLITT-INt 0 X80-LSmitll_SPLITT-OUT-X212-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t992 X80-LSmitll_SPLITT-OUT-X99-LSmitll_DFFT-INt 0 X80-LSmitll_SPLITT-OUT-X99-LSmitll_DFFT-IN 0 z0=5 td=2.7ps
X80 X64-LSmitll_DFFT-OUT-X80-LSmitll_SPLITT-IN X80-LSmitll_SPLITT-OUT-X212-LSmitll_SPLITT-INt X80-LSmitll_SPLITT-OUT-X99-LSmitll_DFFT-INt LSmitll_SPLITT

t993 X81-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-INt 0 X81-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t994 X81-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt 0 X81-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN 0 z0=5 td=2.8ps
X81 X65-LSmitll_AND2T-OUT-X81-LSmitll_SPLITT-IN X81-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-INt X81-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt LSmitll_SPLITT

t995 X82-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt 0 X82-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN 0 z0=5 td=2.8ps
t996 X82-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-INt 0 X82-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
X82 X66-LSmitll_AND2T-OUT-X82-LSmitll_SPLITT-IN X82-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt X82-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-INt LSmitll_SPLITT

t997 X83-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-INt 0 X83-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-IN 0 z0=5 td=1.9ps
t998 X83-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt 0 X83-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN 0 z0=5 td=3.7ps
X83 X67-LSmitll_AND2T-OUT-X83-LSmitll_SPLITT-IN X83-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-INt X83-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt LSmitll_SPLITT

t999 X84-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt 0 X84-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN 0 z0=5 td=4.2ps
t1000 X84-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-INt 0 X84-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
X84 X68-LSmitll_AND2T-OUT-X84-LSmitll_SPLITT-IN X84-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt X84-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-INt LSmitll_SPLITT

t1001 X85-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-INt 0 X85-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-IN 0 z0=5 td=1.4ps
t1002 X85-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-INt 0 X85-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
X85 X69-LSmitll_AND2T-OUT-X85-LSmitll_SPLITT-IN X85-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-INt X85-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-INt LSmitll_SPLITT

t1003 X86-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-INt 0 X86-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-IN 0 z0=5 td=5.3ps
t1004 X86-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt 0 X86-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
X86 X70-LSmitll_AND2T-OUT-X86-LSmitll_SPLITT-IN X86-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-INt X86-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt LSmitll_SPLITT

t1005 X87-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt 0 X87-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN 0 z0=5 td=3.1ps
t1006 X87-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-INt 0 X87-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-IN 0 z0=5 td=4.2ps
X87 X71-LSmitll_AND2T-OUT-X87-LSmitll_SPLITT-IN X87-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt X87-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-INt LSmitll_SPLITT

t1007 X88-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-INt 0 X88-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-IN 0 z0=5 td=3.7ps
t1008 X88-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-INt 0 X88-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-IN 0 z0=5 td=4.0ps
X88 X72-LSmitll_AND2T-OUT-X88-LSmitll_SPLITT-IN X88-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-INt X88-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-INt LSmitll_SPLITT

t1009 X89-LSmitll_DFFT-OUT-X109-LSmitll_SPLITT-INt 0 X89-LSmitll_DFFT-OUT-X109-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X89 X73-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-IN X468-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-IN X89-LSmitll_DFFT-OUT-X109-LSmitll_SPLITT-INt LSmitll_DFFT

t1010 X90-LSmitll_DFFT-OUT-X91-LSmitll_DFFT-INt 0 X90-LSmitll_DFFT-OUT-X91-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X90 X74-LSmitll_SPLITT-OUT-X90-LSmitll_DFFT-IN X468-LSmitll_SPLITT-OUT-X90-LSmitll_DFFT-IN X90-LSmitll_DFFT-OUT-X91-LSmitll_DFFT-INt LSmitll_DFFT

t1011 X91-LSmitll_DFFT-OUT-X110-LSmitll_SPLITT-INt 0 X91-LSmitll_DFFT-OUT-X110-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X91 X90-LSmitll_DFFT-OUT-X91-LSmitll_DFFT-IN X533-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-IN X91-LSmitll_DFFT-OUT-X110-LSmitll_SPLITT-INt LSmitll_DFFT

t1012 X92-LSmitll_DFFT-OUT-X111-LSmitll_SPLITT-INt 0 X92-LSmitll_DFFT-OUT-X111-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
X92 X75-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-IN X461-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-IN X92-LSmitll_DFFT-OUT-X111-LSmitll_SPLITT-INt LSmitll_DFFT

t1013 X93-LSmitll_DFFT-OUT-X94-LSmitll_DFFT-INt 0 X93-LSmitll_DFFT-OUT-X94-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X93 X76-LSmitll_SPLITT-OUT-X93-LSmitll_DFFT-IN X466-LSmitll_SPLITT-OUT-X93-LSmitll_DFFT-IN X93-LSmitll_DFFT-OUT-X94-LSmitll_DFFT-INt LSmitll_DFFT

t1014 X94-LSmitll_DFFT-OUT-X112-LSmitll_SPLITT-INt 0 X94-LSmitll_DFFT-OUT-X112-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X94 X93-LSmitll_DFFT-OUT-X94-LSmitll_DFFT-IN X534-LSmitll_SPLITT-OUT-X94-LSmitll_DFFT-IN X94-LSmitll_DFFT-OUT-X112-LSmitll_SPLITT-INt LSmitll_DFFT

t1015 X95-LSmitll_DFFT-OUT-X113-LSmitll_SPLITT-INt 0 X95-LSmitll_DFFT-OUT-X113-LSmitll_SPLITT-IN 0 z0=5 td=4.6ps
X95 X77-LSmitll_SPLITT-OUT-X95-LSmitll_DFFT-IN X367-LSmitll_SPLITT-OUT-X95-LSmitll_DFFT-IN X95-LSmitll_DFFT-OUT-X113-LSmitll_SPLITT-INt LSmitll_DFFT

t1016 X96-LSmitll_DFFT-OUT-X97-LSmitll_DFFT-INt 0 X96-LSmitll_DFFT-OUT-X97-LSmitll_DFFT-IN 0 z0=5 td=3.9ps
X96 X78-LSmitll_SPLITT-OUT-X96-LSmitll_DFFT-IN X365-LSmitll_SPLITT-OUT-X96-LSmitll_DFFT-IN X96-LSmitll_DFFT-OUT-X97-LSmitll_DFFT-INt LSmitll_DFFT

t1017 X97-LSmitll_DFFT-OUT-X114-LSmitll_SPLITT-INt 0 X97-LSmitll_DFFT-OUT-X114-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X97 X96-LSmitll_DFFT-OUT-X97-LSmitll_DFFT-IN X535-LSmitll_SPLITT-OUT-X97-LSmitll_DFFT-IN X97-LSmitll_DFFT-OUT-X114-LSmitll_SPLITT-INt LSmitll_DFFT

t1018 X98-LSmitll_DFFT-OUT-X115-LSmitll_SPLITT-INt 0 X98-LSmitll_DFFT-OUT-X115-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X98 X79-LSmitll_SPLITT-OUT-X98-LSmitll_DFFT-IN X337-LSmitll_SPLITT-OUT-X98-LSmitll_DFFT-IN X98-LSmitll_DFFT-OUT-X115-LSmitll_SPLITT-INt LSmitll_DFFT

t1019 X99-LSmitll_DFFT-OUT-X100-LSmitll_DFFT-INt 0 X99-LSmitll_DFFT-OUT-X100-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X99 X80-LSmitll_SPLITT-OUT-X99-LSmitll_DFFT-IN X335-LSmitll_SPLITT-OUT-X99-LSmitll_DFFT-IN X99-LSmitll_DFFT-OUT-X100-LSmitll_DFFT-INt LSmitll_DFFT

t1020 X100-LSmitll_DFFT-OUT-X116-LSmitll_SPLITT-INt 0 X100-LSmitll_DFFT-OUT-X116-LSmitll_SPLITT-IN 0 z0=5 td=2.8ps
X100 X99-LSmitll_DFFT-OUT-X100-LSmitll_DFFT-IN X334-LSmitll_SPLITT-OUT-X100-LSmitll_DFFT-IN X100-LSmitll_DFFT-OUT-X116-LSmitll_SPLITT-INt LSmitll_DFFT

t1021 X101-LSmitll_AND2T-OUT-X117-LSmitll_SPLITT-INt 0 X101-LSmitll_AND2T-OUT-X117-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X101 X81-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN X83-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN X359-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN X101-LSmitll_AND2T-OUT-X117-LSmitll_SPLITT-INt LSmitll_AND2T

t1022 X102-LSmitll_AND2T-OUT-X118-LSmitll_SPLITT-INt 0 X102-LSmitll_AND2T-OUT-X118-LSmitll_SPLITT-IN 0 z0=5 td=4.7ps
X102 X81-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-IN X84-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-IN X360-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-IN X102-LSmitll_AND2T-OUT-X118-LSmitll_SPLITT-INt LSmitll_AND2T

t1023 X103-LSmitll_AND2T-OUT-X119-LSmitll_SPLITT-INt 0 X103-LSmitll_AND2T-OUT-X119-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
X103 X83-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-IN X82-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-IN X437-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-IN X103-LSmitll_AND2T-OUT-X119-LSmitll_SPLITT-INt LSmitll_AND2T

t1024 X104-LSmitll_AND2T-OUT-X120-LSmitll_SPLITT-INt 0 X104-LSmitll_AND2T-OUT-X120-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X104 X82-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN X84-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN X442-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN X104-LSmitll_AND2T-OUT-X120-LSmitll_SPLITT-INt LSmitll_AND2T

t1025 X105-LSmitll_AND2T-OUT-X121-LSmitll_SPLITT-INt 0 X105-LSmitll_AND2T-OUT-X121-LSmitll_SPLITT-IN 0 z0=5 td=7.2ps
X105 X85-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-IN X87-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-IN X536-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-IN X105-LSmitll_AND2T-OUT-X121-LSmitll_SPLITT-INt LSmitll_AND2T

t1026 X106-LSmitll_AND2T-OUT-X122-LSmitll_SPLITT-INt 0 X106-LSmitll_AND2T-OUT-X122-LSmitll_SPLITT-IN 0 z0=5 td=7.2ps
X106 X85-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-IN X88-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-IN X537-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-IN X106-LSmitll_AND2T-OUT-X122-LSmitll_SPLITT-INt LSmitll_AND2T

t1027 X107-LSmitll_AND2T-OUT-X123-LSmitll_SPLITT-INt 0 X107-LSmitll_AND2T-OUT-X123-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X107 X87-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN X86-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN X538-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN X107-LSmitll_AND2T-OUT-X123-LSmitll_SPLITT-INt LSmitll_AND2T

t1028 X108-LSmitll_AND2T-OUT-X124-LSmitll_SPLITT-INt 0 X108-LSmitll_AND2T-OUT-X124-LSmitll_SPLITT-IN 0 z0=5 td=7.2ps
X108 X86-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-IN X88-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-IN X412-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-IN X108-LSmitll_AND2T-OUT-X124-LSmitll_SPLITT-INt LSmitll_AND2T

t1029 X109-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-INt 0 X109-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-IN 0 z0=5 td=2.8ps
t1030 X109-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-INt 0 X109-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X109 X89-LSmitll_DFFT-OUT-X109-LSmitll_SPLITT-IN X109-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-INt X109-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-INt LSmitll_SPLITT

t1031 X110-LSmitll_SPLITT-OUT-X192-LSmitll_SPLITT-INt 0 X110-LSmitll_SPLITT-OUT-X192-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
t1032 X110-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-INt 0 X110-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X110 X91-LSmitll_DFFT-OUT-X110-LSmitll_SPLITT-IN X110-LSmitll_SPLITT-OUT-X192-LSmitll_SPLITT-INt X110-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-INt LSmitll_SPLITT

t1033 X111-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt 0 X111-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t1034 X111-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-INt 0 X111-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-IN 0 z0=5 td=8.6ps
X111 X92-LSmitll_DFFT-OUT-X111-LSmitll_SPLITT-IN X111-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt X111-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-INt LSmitll_SPLITT

t1035 X112-LSmitll_SPLITT-OUT-X199-LSmitll_SPLITT-INt 0 X112-LSmitll_SPLITT-OUT-X199-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1036 X112-LSmitll_SPLITT-OUT-X141-LSmitll_DFFT-INt 0 X112-LSmitll_SPLITT-OUT-X141-LSmitll_DFFT-IN 0 z0=5 td=4.0ps
X112 X94-LSmitll_DFFT-OUT-X112-LSmitll_SPLITT-IN X112-LSmitll_SPLITT-OUT-X199-LSmitll_SPLITT-INt X112-LSmitll_SPLITT-OUT-X141-LSmitll_DFFT-INt LSmitll_SPLITT

t1037 X113-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-INt 0 X113-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1038 X113-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-INt 0 X113-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-IN 0 z0=5 td=4.7ps
X113 X95-LSmitll_DFFT-OUT-X113-LSmitll_SPLITT-IN X113-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-INt X113-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-INt LSmitll_SPLITT

t1039 X114-LSmitll_SPLITT-OUT-X206-LSmitll_SPLITT-INt 0 X114-LSmitll_SPLITT-OUT-X206-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1040 X114-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-INt 0 X114-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-IN 0 z0=5 td=2.9ps
X114 X97-LSmitll_DFFT-OUT-X114-LSmitll_SPLITT-IN X114-LSmitll_SPLITT-OUT-X206-LSmitll_SPLITT-INt X114-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-INt LSmitll_SPLITT

t1041 X115-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt 0 X115-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN 0 z0=5 td=3.0ps
t1042 X115-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-INt 0 X115-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-IN 0 z0=5 td=3.6ps
X115 X98-LSmitll_DFFT-OUT-X115-LSmitll_SPLITT-IN X115-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt X115-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-INt LSmitll_SPLITT

t1043 X116-LSmitll_SPLITT-OUT-X213-LSmitll_SPLITT-INt 0 X116-LSmitll_SPLITT-OUT-X213-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
t1044 X116-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-INt 0 X116-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X116 X100-LSmitll_DFFT-OUT-X116-LSmitll_SPLITT-IN X116-LSmitll_SPLITT-OUT-X213-LSmitll_SPLITT-INt X116-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-INt LSmitll_SPLITT

t1045 X117-LSmitll_SPLITT-OUT-X126-LSmitll_SPLITT-INt 0 X117-LSmitll_SPLITT-OUT-X126-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
t1046 X117-LSmitll_SPLITT-OUT-X125-LSmitll_SPLITT-INt 0 X117-LSmitll_SPLITT-OUT-X125-LSmitll_SPLITT-IN 0 z0=5 td=7.6ps
X117 X101-LSmitll_AND2T-OUT-X117-LSmitll_SPLITT-IN X117-LSmitll_SPLITT-OUT-X126-LSmitll_SPLITT-INt X117-LSmitll_SPLITT-OUT-X125-LSmitll_SPLITT-INt LSmitll_SPLITT

t1047 X118-LSmitll_SPLITT-OUT-X283-LSmitll_AND2T-INt 0 X118-LSmitll_SPLITT-OUT-X283-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
t1048 X118-LSmitll_SPLITT-OUT-X127-LSmitll_SPLITT-INt 0 X118-LSmitll_SPLITT-OUT-X127-LSmitll_SPLITT-IN 0 z0=5 td=4.1ps
X118 X102-LSmitll_AND2T-OUT-X118-LSmitll_SPLITT-IN X118-LSmitll_SPLITT-OUT-X283-LSmitll_AND2T-INt X118-LSmitll_SPLITT-OUT-X127-LSmitll_SPLITT-INt LSmitll_SPLITT

t1049 X119-LSmitll_SPLITT-OUT-X129-LSmitll_SPLITT-INt 0 X119-LSmitll_SPLITT-OUT-X129-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1050 X119-LSmitll_SPLITT-OUT-X128-LSmitll_SPLITT-INt 0 X119-LSmitll_SPLITT-OUT-X128-LSmitll_SPLITT-IN 0 z0=5 td=6.8ps
X119 X103-LSmitll_AND2T-OUT-X119-LSmitll_SPLITT-IN X119-LSmitll_SPLITT-OUT-X129-LSmitll_SPLITT-INt X119-LSmitll_SPLITT-OUT-X128-LSmitll_SPLITT-INt LSmitll_SPLITT

t1051 X120-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-INt 0 X120-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1052 X120-LSmitll_SPLITT-OUT-X130-LSmitll_SPLITT-INt 0 X120-LSmitll_SPLITT-OUT-X130-LSmitll_SPLITT-IN 0 z0=5 td=4.3ps
X120 X104-LSmitll_AND2T-OUT-X120-LSmitll_SPLITT-IN X120-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-INt X120-LSmitll_SPLITT-OUT-X130-LSmitll_SPLITT-INt LSmitll_SPLITT

t1053 X121-LSmitll_SPLITT-OUT-X300-LSmitll_AND2T-INt 0 X121-LSmitll_SPLITT-OUT-X300-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1054 X121-LSmitll_SPLITT-OUT-X131-LSmitll_SPLITT-INt 0 X121-LSmitll_SPLITT-OUT-X131-LSmitll_SPLITT-IN 0 z0=5 td=3.4ps
X121 X105-LSmitll_AND2T-OUT-X121-LSmitll_SPLITT-IN X121-LSmitll_SPLITT-OUT-X300-LSmitll_AND2T-INt X121-LSmitll_SPLITT-OUT-X131-LSmitll_SPLITT-INt LSmitll_SPLITT

t1055 X122-LSmitll_SPLITT-OUT-X133-LSmitll_SPLITT-INt 0 X122-LSmitll_SPLITT-OUT-X133-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1056 X122-LSmitll_SPLITT-OUT-X132-LSmitll_SPLITT-INt 0 X122-LSmitll_SPLITT-OUT-X132-LSmitll_SPLITT-IN 0 z0=5 td=6.0ps
X122 X106-LSmitll_AND2T-OUT-X122-LSmitll_SPLITT-IN X122-LSmitll_SPLITT-OUT-X133-LSmitll_SPLITT-INt X122-LSmitll_SPLITT-OUT-X132-LSmitll_SPLITT-INt LSmitll_SPLITT

t1057 X123-LSmitll_SPLITT-OUT-X298-LSmitll_AND2T-INt 0 X123-LSmitll_SPLITT-OUT-X298-LSmitll_AND2T-IN 0 z0=5 td=8.0ps
t1058 X123-LSmitll_SPLITT-OUT-X134-LSmitll_SPLITT-INt 0 X123-LSmitll_SPLITT-OUT-X134-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X123 X107-LSmitll_AND2T-OUT-X123-LSmitll_SPLITT-IN X123-LSmitll_SPLITT-OUT-X298-LSmitll_AND2T-INt X123-LSmitll_SPLITT-OUT-X134-LSmitll_SPLITT-INt LSmitll_SPLITT

t1059 X124-LSmitll_SPLITT-OUT-X136-LSmitll_SPLITT-INt 0 X124-LSmitll_SPLITT-OUT-X136-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1060 X124-LSmitll_SPLITT-OUT-X135-LSmitll_SPLITT-INt 0 X124-LSmitll_SPLITT-OUT-X135-LSmitll_SPLITT-IN 0 z0=5 td=19.2ps
X124 X108-LSmitll_AND2T-OUT-X124-LSmitll_SPLITT-IN X124-LSmitll_SPLITT-OUT-X136-LSmitll_SPLITT-INt X124-LSmitll_SPLITT-OUT-X135-LSmitll_SPLITT-INt LSmitll_SPLITT

t1061 X125-LSmitll_SPLITT-OUT-X280-LSmitll_AND2T-INt 0 X125-LSmitll_SPLITT-OUT-X280-LSmitll_AND2T-IN 0 z0=5 td=3.9ps
t1062 X125-LSmitll_SPLITT-OUT-X276-LSmitll_AND2T-INt 0 X125-LSmitll_SPLITT-OUT-X276-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
X125 X117-LSmitll_SPLITT-OUT-X125-LSmitll_SPLITT-IN X125-LSmitll_SPLITT-OUT-X280-LSmitll_AND2T-INt X125-LSmitll_SPLITT-OUT-X276-LSmitll_AND2T-INt LSmitll_SPLITT

t1063 X126-LSmitll_SPLITT-OUT-X288-LSmitll_AND2T-INt 0 X126-LSmitll_SPLITT-OUT-X288-LSmitll_AND2T-IN 0 z0=5 td=3.8ps
t1064 X126-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-INt 0 X126-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X126 X117-LSmitll_SPLITT-OUT-X126-LSmitll_SPLITT-IN X126-LSmitll_SPLITT-OUT-X288-LSmitll_AND2T-INt X126-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-INt LSmitll_SPLITT

t1065 X127-LSmitll_SPLITT-OUT-X279-LSmitll_AND2T-INt 0 X127-LSmitll_SPLITT-OUT-X279-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1066 X127-LSmitll_SPLITT-OUT-X275-LSmitll_AND2T-INt 0 X127-LSmitll_SPLITT-OUT-X275-LSmitll_AND2T-IN 0 z0=5 td=5.4ps
X127 X118-LSmitll_SPLITT-OUT-X127-LSmitll_SPLITT-IN X127-LSmitll_SPLITT-OUT-X279-LSmitll_AND2T-INt X127-LSmitll_SPLITT-OUT-X275-LSmitll_AND2T-INt LSmitll_SPLITT

t1067 X128-LSmitll_SPLITT-OUT-X278-LSmitll_AND2T-INt 0 X128-LSmitll_SPLITT-OUT-X278-LSmitll_AND2T-IN 0 z0=5 td=4.3ps
t1068 X128-LSmitll_SPLITT-OUT-X274-LSmitll_AND2T-INt 0 X128-LSmitll_SPLITT-OUT-X274-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
X128 X119-LSmitll_SPLITT-OUT-X128-LSmitll_SPLITT-IN X128-LSmitll_SPLITT-OUT-X278-LSmitll_AND2T-INt X128-LSmitll_SPLITT-OUT-X274-LSmitll_AND2T-INt LSmitll_SPLITT

t1069 X129-LSmitll_SPLITT-OUT-X286-LSmitll_AND2T-INt 0 X129-LSmitll_SPLITT-OUT-X286-LSmitll_AND2T-IN 0 z0=5 td=4.6ps
t1070 X129-LSmitll_SPLITT-OUT-X282-LSmitll_AND2T-INt 0 X129-LSmitll_SPLITT-OUT-X282-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X129 X119-LSmitll_SPLITT-OUT-X129-LSmitll_SPLITT-IN X129-LSmitll_SPLITT-OUT-X286-LSmitll_AND2T-INt X129-LSmitll_SPLITT-OUT-X282-LSmitll_AND2T-INt LSmitll_SPLITT

t1071 X130-LSmitll_SPLITT-OUT-X277-LSmitll_AND2T-INt 0 X130-LSmitll_SPLITT-OUT-X277-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t1072 X130-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-INt 0 X130-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-IN 0 z0=5 td=3.8ps
X130 X120-LSmitll_SPLITT-OUT-X130-LSmitll_SPLITT-IN X130-LSmitll_SPLITT-OUT-X277-LSmitll_AND2T-INt X130-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-INt LSmitll_SPLITT

t1073 X131-LSmitll_SPLITT-OUT-X296-LSmitll_AND2T-INt 0 X131-LSmitll_SPLITT-OUT-X296-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1074 X131-LSmitll_SPLITT-OUT-X292-LSmitll_AND2T-INt 0 X131-LSmitll_SPLITT-OUT-X292-LSmitll_AND2T-IN 0 z0=5 td=3.4ps
X131 X121-LSmitll_SPLITT-OUT-X131-LSmitll_SPLITT-IN X131-LSmitll_SPLITT-OUT-X296-LSmitll_AND2T-INt X131-LSmitll_SPLITT-OUT-X292-LSmitll_AND2T-INt LSmitll_SPLITT

t1075 X132-LSmitll_SPLITT-OUT-X291-LSmitll_AND2T-INt 0 X132-LSmitll_SPLITT-OUT-X291-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1076 X132-LSmitll_SPLITT-OUT-X287-LSmitll_AND2T-INt 0 X132-LSmitll_SPLITT-OUT-X287-LSmitll_AND2T-IN 0 z0=5 td=4.9ps
X132 X122-LSmitll_SPLITT-OUT-X132-LSmitll_SPLITT-IN X132-LSmitll_SPLITT-OUT-X291-LSmitll_AND2T-INt X132-LSmitll_SPLITT-OUT-X287-LSmitll_AND2T-INt LSmitll_SPLITT

t1077 X133-LSmitll_SPLITT-OUT-X299-LSmitll_AND2T-INt 0 X133-LSmitll_SPLITT-OUT-X299-LSmitll_AND2T-IN 0 z0=5 td=9.4ps
t1078 X133-LSmitll_SPLITT-OUT-X295-LSmitll_AND2T-INt 0 X133-LSmitll_SPLITT-OUT-X295-LSmitll_AND2T-IN 0 z0=5 td=3.2ps
X133 X122-LSmitll_SPLITT-OUT-X133-LSmitll_SPLITT-IN X133-LSmitll_SPLITT-OUT-X299-LSmitll_AND2T-INt X133-LSmitll_SPLITT-OUT-X295-LSmitll_AND2T-INt LSmitll_SPLITT

t1079 X134-LSmitll_SPLITT-OUT-X294-LSmitll_AND2T-INt 0 X134-LSmitll_SPLITT-OUT-X294-LSmitll_AND2T-IN 0 z0=5 td=4.6ps
t1080 X134-LSmitll_SPLITT-OUT-X290-LSmitll_AND2T-INt 0 X134-LSmitll_SPLITT-OUT-X290-LSmitll_AND2T-IN 0 z0=5 td=2.9ps
X134 X123-LSmitll_SPLITT-OUT-X134-LSmitll_SPLITT-IN X134-LSmitll_SPLITT-OUT-X294-LSmitll_AND2T-INt X134-LSmitll_SPLITT-OUT-X290-LSmitll_AND2T-INt LSmitll_SPLITT

t1081 X135-LSmitll_SPLITT-OUT-X289-LSmitll_AND2T-INt 0 X135-LSmitll_SPLITT-OUT-X289-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t1082 X135-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-INt 0 X135-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-IN 0 z0=5 td=4.5ps
X135 X124-LSmitll_SPLITT-OUT-X135-LSmitll_SPLITT-IN X135-LSmitll_SPLITT-OUT-X289-LSmitll_AND2T-INt X135-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-INt LSmitll_SPLITT

t1083 X136-LSmitll_SPLITT-OUT-X297-LSmitll_AND2T-INt 0 X136-LSmitll_SPLITT-OUT-X297-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1084 X136-LSmitll_SPLITT-OUT-X293-LSmitll_AND2T-INt 0 X136-LSmitll_SPLITT-OUT-X293-LSmitll_AND2T-IN 0 z0=5 td=7.1ps
X136 X124-LSmitll_SPLITT-OUT-X136-LSmitll_SPLITT-IN X136-LSmitll_SPLITT-OUT-X297-LSmitll_AND2T-INt X136-LSmitll_SPLITT-OUT-X293-LSmitll_AND2T-INt LSmitll_SPLITT

t1085 X137-LSmitll_DFFT-OUT-X149-LSmitll_SPLITT-INt 0 X137-LSmitll_DFFT-OUT-X149-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X137 X109-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-IN X539-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-IN X137-LSmitll_DFFT-OUT-X149-LSmitll_SPLITT-INt LSmitll_DFFT

t1086 X138-LSmitll_DFFT-OUT-X139-LSmitll_DFFT-INt 0 X138-LSmitll_DFFT-OUT-X139-LSmitll_DFFT-IN 0 z0=5 td=2.4ps
X138 X110-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-IN X505-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-IN X138-LSmitll_DFFT-OUT-X139-LSmitll_DFFT-INt LSmitll_DFFT

t1087 X139-LSmitll_DFFT-OUT-X150-LSmitll_SPLITT-INt 0 X139-LSmitll_DFFT-OUT-X150-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X139 X138-LSmitll_DFFT-OUT-X139-LSmitll_DFFT-IN X540-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-IN X139-LSmitll_DFFT-OUT-X150-LSmitll_SPLITT-INt LSmitll_DFFT

t1088 X140-LSmitll_DFFT-OUT-X151-LSmitll_SPLITT-INt 0 X140-LSmitll_DFFT-OUT-X151-LSmitll_SPLITT-IN 0 z0=5 td=8.8ps
X140 X111-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-IN X474-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-IN X140-LSmitll_DFFT-OUT-X151-LSmitll_SPLITT-INt LSmitll_DFFT

t1089 X141-LSmitll_DFFT-OUT-X142-LSmitll_DFFT-INt 0 X141-LSmitll_DFFT-OUT-X142-LSmitll_DFFT-IN 0 z0=5 td=6.7ps
X141 X112-LSmitll_SPLITT-OUT-X141-LSmitll_DFFT-IN X439-LSmitll_SPLITT-OUT-X141-LSmitll_DFFT-IN X141-LSmitll_DFFT-OUT-X142-LSmitll_DFFT-INt LSmitll_DFFT

t1090 X142-LSmitll_DFFT-OUT-X152-LSmitll_SPLITT-INt 0 X142-LSmitll_DFFT-OUT-X152-LSmitll_SPLITT-IN 0 z0=5 td=28.2ps
X142 X141-LSmitll_DFFT-OUT-X142-LSmitll_DFFT-IN X541-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-IN X142-LSmitll_DFFT-OUT-X152-LSmitll_SPLITT-INt LSmitll_DFFT

t1091 X143-LSmitll_DFFT-OUT-X153-LSmitll_SPLITT-INt 0 X143-LSmitll_DFFT-OUT-X153-LSmitll_SPLITT-IN 0 z0=5 td=6.6ps
X143 X113-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-IN X404-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-IN X143-LSmitll_DFFT-OUT-X153-LSmitll_SPLITT-INt LSmitll_DFFT

t1092 X144-LSmitll_DFFT-OUT-X145-LSmitll_DFFT-INt 0 X144-LSmitll_DFFT-OUT-X145-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X144 X114-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-IN X398-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-IN X144-LSmitll_DFFT-OUT-X145-LSmitll_DFFT-INt LSmitll_DFFT

t1093 X145-LSmitll_DFFT-OUT-X154-LSmitll_SPLITT-INt 0 X145-LSmitll_DFFT-OUT-X154-LSmitll_SPLITT-IN 0 z0=5 td=7.3ps
X145 X144-LSmitll_DFFT-OUT-X145-LSmitll_DFFT-IN X399-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-IN X145-LSmitll_DFFT-OUT-X154-LSmitll_SPLITT-INt LSmitll_DFFT

t1094 X146-LSmitll_DFFT-OUT-X155-LSmitll_SPLITT-INt 0 X146-LSmitll_DFFT-OUT-X155-LSmitll_SPLITT-IN 0 z0=5 td=6.4ps
X146 X115-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-IN X373-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-IN X146-LSmitll_DFFT-OUT-X155-LSmitll_SPLITT-INt LSmitll_DFFT

t1095 X147-LSmitll_DFFT-OUT-X148-LSmitll_DFFT-INt 0 X147-LSmitll_DFFT-OUT-X148-LSmitll_DFFT-IN 0 z0=5 td=3.6ps
X147 X116-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-IN X337-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-IN X147-LSmitll_DFFT-OUT-X148-LSmitll_DFFT-INt LSmitll_DFFT

t1096 X148-LSmitll_DFFT-OUT-X156-LSmitll_SPLITT-INt 0 X148-LSmitll_DFFT-OUT-X156-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
X148 X147-LSmitll_DFFT-OUT-X148-LSmitll_DFFT-IN X373-LSmitll_SPLITT-OUT-X148-LSmitll_DFFT-IN X148-LSmitll_DFFT-OUT-X156-LSmitll_SPLITT-INt LSmitll_DFFT

t1097 X149-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-INt 0 X149-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t1098 X149-LSmitll_SPLITT-OUT-X157-LSmitll_DFFT-INt 0 X149-LSmitll_SPLITT-OUT-X157-LSmitll_DFFT-IN 0 z0=5 td=2.8ps
X149 X137-LSmitll_DFFT-OUT-X149-LSmitll_SPLITT-IN X149-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-INt X149-LSmitll_SPLITT-OUT-X157-LSmitll_DFFT-INt LSmitll_SPLITT

t1099 X150-LSmitll_SPLITT-OUT-X193-LSmitll_SPLITT-INt 0 X150-LSmitll_SPLITT-OUT-X193-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
t1100 X150-LSmitll_SPLITT-OUT-X158-LSmitll_DFFT-INt 0 X150-LSmitll_SPLITT-OUT-X158-LSmitll_DFFT-IN 0 z0=5 td=3.5ps
X150 X139-LSmitll_DFFT-OUT-X150-LSmitll_SPLITT-IN X150-LSmitll_SPLITT-OUT-X193-LSmitll_SPLITT-INt X150-LSmitll_SPLITT-OUT-X158-LSmitll_DFFT-INt LSmitll_SPLITT

t1101 X151-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt 0 X151-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
t1102 X151-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-INt 0 X151-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-IN 0 z0=5 td=4.0ps
X151 X140-LSmitll_DFFT-OUT-X151-LSmitll_SPLITT-IN X151-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt X151-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-INt LSmitll_SPLITT

t1103 X152-LSmitll_SPLITT-OUT-X200-LSmitll_SPLITT-INt 0 X152-LSmitll_SPLITT-OUT-X200-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1104 X152-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-INt 0 X152-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X152 X142-LSmitll_DFFT-OUT-X152-LSmitll_SPLITT-IN X152-LSmitll_SPLITT-OUT-X200-LSmitll_SPLITT-INt X152-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-INt LSmitll_SPLITT

t1105 X153-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-INt 0 X153-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1106 X153-LSmitll_SPLITT-OUT-X163-LSmitll_DFFT-INt 0 X153-LSmitll_SPLITT-OUT-X163-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X153 X143-LSmitll_DFFT-OUT-X153-LSmitll_SPLITT-IN X153-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-INt X153-LSmitll_SPLITT-OUT-X163-LSmitll_DFFT-INt LSmitll_SPLITT

t1107 X154-LSmitll_SPLITT-OUT-X207-LSmitll_SPLITT-INt 0 X154-LSmitll_SPLITT-OUT-X207-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1108 X154-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-INt 0 X154-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-IN 0 z0=5 td=6.2ps
X154 X145-LSmitll_DFFT-OUT-X154-LSmitll_SPLITT-IN X154-LSmitll_SPLITT-OUT-X207-LSmitll_SPLITT-INt X154-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-INt LSmitll_SPLITT

t1109 X155-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-INt 0 X155-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-IN 0 z0=5 td=13.2ps
t1110 X155-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-INt 0 X155-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-IN 0 z0=5 td=3.0ps
X155 X146-LSmitll_DFFT-OUT-X155-LSmitll_SPLITT-IN X155-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-INt X155-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-INt LSmitll_SPLITT

t1111 X156-LSmitll_SPLITT-OUT-X214-LSmitll_SPLITT-INt 0 X156-LSmitll_SPLITT-OUT-X214-LSmitll_SPLITT-IN 0 z0=5 td=4.6ps
t1112 X156-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-INt 0 X156-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X156 X148-LSmitll_DFFT-OUT-X156-LSmitll_SPLITT-IN X156-LSmitll_SPLITT-OUT-X214-LSmitll_SPLITT-INt X156-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-INt LSmitll_SPLITT

t1113 X157-LSmitll_DFFT-OUT-X169-LSmitll_SPLITT-INt 0 X157-LSmitll_DFFT-OUT-X169-LSmitll_SPLITT-IN 0 z0=5 td=3.5ps
X157 X149-LSmitll_SPLITT-OUT-X157-LSmitll_DFFT-IN X507-LSmitll_SPLITT-OUT-X157-LSmitll_DFFT-IN X157-LSmitll_DFFT-OUT-X169-LSmitll_SPLITT-INt LSmitll_DFFT

t1114 X158-LSmitll_DFFT-OUT-X159-LSmitll_DFFT-INt 0 X158-LSmitll_DFFT-OUT-X159-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X158 X150-LSmitll_SPLITT-OUT-X158-LSmitll_DFFT-IN X507-LSmitll_SPLITT-OUT-X158-LSmitll_DFFT-IN X158-LSmitll_DFFT-OUT-X159-LSmitll_DFFT-INt LSmitll_DFFT

t1115 X159-LSmitll_DFFT-OUT-X170-LSmitll_SPLITT-INt 0 X159-LSmitll_DFFT-OUT-X170-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X159 X158-LSmitll_DFFT-OUT-X159-LSmitll_DFFT-IN X542-LSmitll_SPLITT-OUT-X159-LSmitll_DFFT-IN X159-LSmitll_DFFT-OUT-X170-LSmitll_SPLITT-INt LSmitll_DFFT

t1116 X160-LSmitll_DFFT-OUT-X171-LSmitll_SPLITT-INt 0 X160-LSmitll_DFFT-OUT-X171-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X160 X151-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-IN X513-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-IN X160-LSmitll_DFFT-OUT-X171-LSmitll_SPLITT-INt LSmitll_DFFT

t1117 X161-LSmitll_DFFT-OUT-X162-LSmitll_DFFT-INt 0 X161-LSmitll_DFFT-OUT-X162-LSmitll_DFFT-IN 0 z0=5 td=4.0ps
X161 X152-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-IN X385-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-IN X161-LSmitll_DFFT-OUT-X162-LSmitll_DFFT-INt LSmitll_DFFT

t1118 X162-LSmitll_DFFT-OUT-X172-LSmitll_SPLITT-INt 0 X162-LSmitll_DFFT-OUT-X172-LSmitll_SPLITT-IN 0 z0=5 td=13.1ps
X162 X161-LSmitll_DFFT-OUT-X162-LSmitll_DFFT-IN X388-LSmitll_SPLITT-OUT-X162-LSmitll_DFFT-IN X162-LSmitll_DFFT-OUT-X172-LSmitll_SPLITT-INt LSmitll_DFFT

t1119 X163-LSmitll_DFFT-OUT-X173-LSmitll_SPLITT-INt 0 X163-LSmitll_DFFT-OUT-X173-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X163 X153-LSmitll_SPLITT-OUT-X163-LSmitll_DFFT-IN X480-LSmitll_SPLITT-OUT-X163-LSmitll_DFFT-IN X163-LSmitll_DFFT-OUT-X173-LSmitll_SPLITT-INt LSmitll_DFFT

t1120 X164-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-INt 0 X164-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X164 X154-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-IN X482-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-IN X164-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-INt LSmitll_DFFT

t1121 X165-LSmitll_DFFT-OUT-X174-LSmitll_SPLITT-INt 0 X165-LSmitll_DFFT-OUT-X174-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X165 X164-LSmitll_DFFT-OUT-X165-LSmitll_DFFT-IN X543-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-IN X165-LSmitll_DFFT-OUT-X174-LSmitll_SPLITT-INt LSmitll_DFFT

t1122 X166-LSmitll_DFFT-OUT-X175-LSmitll_SPLITT-INt 0 X166-LSmitll_DFFT-OUT-X175-LSmitll_SPLITT-IN 0 z0=5 td=4.0ps
X166 X155-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-IN X544-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-IN X166-LSmitll_DFFT-OUT-X175-LSmitll_SPLITT-INt LSmitll_DFFT

t1123 X167-LSmitll_DFFT-OUT-X168-LSmitll_DFFT-INt 0 X167-LSmitll_DFFT-OUT-X168-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X167 X156-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-IN X374-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-IN X167-LSmitll_DFFT-OUT-X168-LSmitll_DFFT-INt LSmitll_DFFT

t1124 X168-LSmitll_DFFT-OUT-X176-LSmitll_SPLITT-INt 0 X168-LSmitll_DFFT-OUT-X176-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
X168 X167-LSmitll_DFFT-OUT-X168-LSmitll_DFFT-IN X379-LSmitll_SPLITT-OUT-X168-LSmitll_DFFT-IN X168-LSmitll_DFFT-OUT-X176-LSmitll_SPLITT-INt LSmitll_DFFT

t1125 X169-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-INt 0 X169-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
t1126 X169-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-INt 0 X169-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-IN 0 z0=5 td=2.9ps
X169 X157-LSmitll_DFFT-OUT-X169-LSmitll_SPLITT-IN X169-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-INt X169-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-INt LSmitll_SPLITT

t1127 X170-LSmitll_SPLITT-OUT-X194-LSmitll_SPLITT-INt 0 X170-LSmitll_SPLITT-OUT-X194-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1128 X170-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-INt 0 X170-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-IN 0 z0=5 td=5.5ps
X170 X159-LSmitll_DFFT-OUT-X170-LSmitll_SPLITT-IN X170-LSmitll_SPLITT-OUT-X194-LSmitll_SPLITT-INt X170-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-INt LSmitll_SPLITT

t1129 X171-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-INt 0 X171-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t1130 X171-LSmitll_SPLITT-OUT-X180-LSmitll_DFFT-INt 0 X171-LSmitll_SPLITT-OUT-X180-LSmitll_DFFT-IN 0 z0=5 td=2.4ps
X171 X160-LSmitll_DFFT-OUT-X171-LSmitll_SPLITT-IN X171-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-INt X171-LSmitll_SPLITT-OUT-X180-LSmitll_DFFT-INt LSmitll_SPLITT

t1131 X172-LSmitll_SPLITT-OUT-X201-LSmitll_SPLITT-INt 0 X172-LSmitll_SPLITT-OUT-X201-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
t1132 X172-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-INt 0 X172-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
X172 X162-LSmitll_DFFT-OUT-X172-LSmitll_SPLITT-IN X172-LSmitll_SPLITT-OUT-X201-LSmitll_SPLITT-INt X172-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-INt LSmitll_SPLITT

t1133 X173-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-INt 0 X173-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
t1134 X173-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-INt 0 X173-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-IN 0 z0=5 td=5.9ps
X173 X163-LSmitll_DFFT-OUT-X173-LSmitll_SPLITT-IN X173-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-INt X173-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-INt LSmitll_SPLITT

t1135 X174-LSmitll_SPLITT-OUT-X208-LSmitll_SPLITT-INt 0 X174-LSmitll_SPLITT-OUT-X208-LSmitll_SPLITT-IN 0 z0=5 td=4.7ps
t1136 X174-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-INt 0 X174-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-IN 0 z0=5 td=3.8ps
X174 X165-LSmitll_DFFT-OUT-X174-LSmitll_SPLITT-IN X174-LSmitll_SPLITT-OUT-X208-LSmitll_SPLITT-INt X174-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-INt LSmitll_SPLITT

t1137 X175-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-INt 0 X175-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-IN 0 z0=5 td=1.7ps
t1138 X175-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-INt 0 X175-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X175 X166-LSmitll_DFFT-OUT-X175-LSmitll_SPLITT-IN X175-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-INt X175-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-INt LSmitll_SPLITT

t1139 X176-LSmitll_SPLITT-OUT-X215-LSmitll_SPLITT-INt 0 X176-LSmitll_SPLITT-OUT-X215-LSmitll_SPLITT-IN 0 z0=5 td=5.9ps
t1140 X176-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-INt 0 X176-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X176 X168-LSmitll_DFFT-OUT-X176-LSmitll_SPLITT-IN X176-LSmitll_SPLITT-OUT-X215-LSmitll_SPLITT-INt X176-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-INt LSmitll_SPLITT

t1141 X177-LSmitll_DFFT-OUT-X230-LSmitll_AND2T-INt 0 X177-LSmitll_DFFT-OUT-X230-LSmitll_AND2T-IN 0 z0=5 td=3.8ps
X177 X169-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-IN X511-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-IN X177-LSmitll_DFFT-OUT-X230-LSmitll_AND2T-INt LSmitll_DFFT

t1142 X178-LSmitll_DFFT-OUT-X179-LSmitll_DFFT-INt 0 X178-LSmitll_DFFT-OUT-X179-LSmitll_DFFT-IN 0 z0=5 td=2.5ps
X178 X170-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-IN X511-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-IN X178-LSmitll_DFFT-OUT-X179-LSmitll_DFFT-INt LSmitll_DFFT

t1143 X179-LSmitll_DFFT-OUT-X195-LSmitll_SPLITT-INt 0 X179-LSmitll_DFFT-OUT-X195-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X179 X178-LSmitll_DFFT-OUT-X179-LSmitll_DFFT-IN X545-LSmitll_SPLITT-OUT-X179-LSmitll_DFFT-IN X179-LSmitll_DFFT-OUT-X195-LSmitll_SPLITT-INt LSmitll_DFFT

t1144 X180-LSmitll_DFFT-OUT-X244-LSmitll_AND2T-INt 0 X180-LSmitll_DFFT-OUT-X244-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X180 X171-LSmitll_SPLITT-OUT-X180-LSmitll_DFFT-IN X546-LSmitll_SPLITT-OUT-X180-LSmitll_DFFT-IN X180-LSmitll_DFFT-OUT-X244-LSmitll_AND2T-INt LSmitll_DFFT

t1145 X181-LSmitll_DFFT-OUT-X182-LSmitll_DFFT-INt 0 X181-LSmitll_DFFT-OUT-X182-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X181 X172-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-IN X417-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-IN X181-LSmitll_DFFT-OUT-X182-LSmitll_DFFT-INt LSmitll_DFFT

t1146 X182-LSmitll_DFFT-OUT-X202-LSmitll_SPLITT-INt 0 X182-LSmitll_DFFT-OUT-X202-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
X182 X181-LSmitll_DFFT-OUT-X182-LSmitll_DFFT-IN X417-LSmitll_SPLITT-OUT-X182-LSmitll_DFFT-IN X182-LSmitll_DFFT-OUT-X202-LSmitll_SPLITT-INt LSmitll_DFFT

t1147 X183-LSmitll_DFFT-OUT-X258-LSmitll_AND2T-INt 0 X183-LSmitll_DFFT-OUT-X258-LSmitll_AND2T-IN 0 z0=5 td=4.5ps
X183 X173-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-IN X500-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-IN X183-LSmitll_DFFT-OUT-X258-LSmitll_AND2T-INt LSmitll_DFFT

t1148 X184-LSmitll_DFFT-OUT-X185-LSmitll_DFFT-INt 0 X184-LSmitll_DFFT-OUT-X185-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X184 X174-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-IN X502-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-IN X184-LSmitll_DFFT-OUT-X185-LSmitll_DFFT-INt LSmitll_DFFT

t1149 X185-LSmitll_DFFT-OUT-X209-LSmitll_SPLITT-INt 0 X185-LSmitll_DFFT-OUT-X209-LSmitll_SPLITT-IN 0 z0=5 td=4.8ps
X185 X184-LSmitll_DFFT-OUT-X185-LSmitll_DFFT-IN X505-LSmitll_SPLITT-OUT-X185-LSmitll_DFFT-IN X185-LSmitll_DFFT-OUT-X209-LSmitll_SPLITT-INt LSmitll_DFFT

t1150 X186-LSmitll_DFFT-OUT-X272-LSmitll_AND2T-INt 0 X186-LSmitll_DFFT-OUT-X272-LSmitll_AND2T-IN 0 z0=5 td=4.8ps
X186 X175-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-IN X376-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-IN X186-LSmitll_DFFT-OUT-X272-LSmitll_AND2T-INt LSmitll_DFFT

t1151 X187-LSmitll_DFFT-OUT-X188-LSmitll_DFFT-INt 0 X187-LSmitll_DFFT-OUT-X188-LSmitll_DFFT-IN 0 z0=5 td=3.8ps
X187 X176-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-IN X376-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-IN X187-LSmitll_DFFT-OUT-X188-LSmitll_DFFT-INt LSmitll_DFFT

t1152 X188-LSmitll_DFFT-OUT-X216-LSmitll_SPLITT-INt 0 X188-LSmitll_DFFT-OUT-X216-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
X188 X187-LSmitll_DFFT-OUT-X188-LSmitll_DFFT-IN X385-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-IN X188-LSmitll_DFFT-OUT-X216-LSmitll_SPLITT-INt LSmitll_DFFT

t1153 X189-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-INt 0 X189-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-IN 0 z0=5 td=1.4ps
t1154 X189-LSmitll_SPLITT-OUT-X217-LSmitll_NDROT-INt 0 X189-LSmitll_SPLITT-OUT-X217-LSmitll_NDROT-IN 0 z0=5 td=2.8ps
X189 X1-LSmitll_SPLITT-OUT-X189-LSmitll_SPLITT-IN X189-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-INt X189-LSmitll_SPLITT-OUT-X217-LSmitll_NDROT-INt LSmitll_SPLITT

t1155 X190-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-INt 0 X190-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t1156 X190-LSmitll_SPLITT-OUT-X219-LSmitll_NDROT-INt 0 X190-LSmitll_SPLITT-OUT-X219-LSmitll_NDROT-IN 0 z0=5 td=2.6ps
X190 X42-LSmitll_SPLITT-OUT-X190-LSmitll_SPLITT-IN X190-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-INt X190-LSmitll_SPLITT-OUT-X219-LSmitll_NDROT-INt LSmitll_SPLITT

t1157 X191-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-INt 0 X191-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t1158 X191-LSmitll_SPLITT-OUT-X221-LSmitll_NDROT-INt 0 X191-LSmitll_SPLITT-OUT-X221-LSmitll_NDROT-IN 0 z0=5 td=2.6ps
X191 X74-LSmitll_SPLITT-OUT-X191-LSmitll_SPLITT-IN X191-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-INt X191-LSmitll_SPLITT-OUT-X221-LSmitll_NDROT-INt LSmitll_SPLITT

t1159 X192-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-INt 0 X192-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1160 X192-LSmitll_SPLITT-OUT-X223-LSmitll_NDROT-INt 0 X192-LSmitll_SPLITT-OUT-X223-LSmitll_NDROT-IN 0 z0=5 td=1.0ps
X192 X110-LSmitll_SPLITT-OUT-X192-LSmitll_SPLITT-IN X192-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-INt X192-LSmitll_SPLITT-OUT-X223-LSmitll_NDROT-INt LSmitll_SPLITT

t1161 X193-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-INt 0 X193-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
t1162 X193-LSmitll_SPLITT-OUT-X225-LSmitll_NDROT-INt 0 X193-LSmitll_SPLITT-OUT-X225-LSmitll_NDROT-IN 0 z0=5 td=2.6ps
X193 X150-LSmitll_SPLITT-OUT-X193-LSmitll_SPLITT-IN X193-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-INt X193-LSmitll_SPLITT-OUT-X225-LSmitll_NDROT-INt LSmitll_SPLITT

t1163 X194-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-INt 0 X194-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t1164 X194-LSmitll_SPLITT-OUT-X227-LSmitll_NDROT-INt 0 X194-LSmitll_SPLITT-OUT-X227-LSmitll_NDROT-IN 0 z0=5 td=2.6ps
X194 X170-LSmitll_SPLITT-OUT-X194-LSmitll_SPLITT-IN X194-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-INt X194-LSmitll_SPLITT-OUT-X227-LSmitll_NDROT-INt LSmitll_SPLITT

t1165 X195-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-INt 0 X195-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t1166 X195-LSmitll_SPLITT-OUT-X229-LSmitll_NDROT-INt 0 X195-LSmitll_SPLITT-OUT-X229-LSmitll_NDROT-IN 0 z0=5 td=2.6ps
X195 X179-LSmitll_DFFT-OUT-X195-LSmitll_SPLITT-IN X195-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-INt X195-LSmitll_SPLITT-OUT-X229-LSmitll_NDROT-INt LSmitll_SPLITT

t1167 X196-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-INt 0 X196-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t1168 X196-LSmitll_SPLITT-OUT-X231-LSmitll_NDROT-INt 0 X196-LSmitll_SPLITT-OUT-X231-LSmitll_NDROT-IN 0 z0=5 td=3.7ps
X196 X3-LSmitll_SPLITT-OUT-X196-LSmitll_SPLITT-IN X196-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-INt X196-LSmitll_SPLITT-OUT-X231-LSmitll_NDROT-INt LSmitll_SPLITT

t1169 X197-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt 0 X197-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN 0 z0=5 td=1.4ps
t1170 X197-LSmitll_SPLITT-OUT-X233-LSmitll_NDROT-INt 0 X197-LSmitll_SPLITT-OUT-X233-LSmitll_NDROT-IN 0 z0=5 td=2.1ps
X197 X44-LSmitll_SPLITT-OUT-X197-LSmitll_SPLITT-IN X197-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt X197-LSmitll_SPLITT-OUT-X233-LSmitll_NDROT-INt LSmitll_SPLITT

t1171 X198-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-INt 0 X198-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
t1172 X198-LSmitll_SPLITT-OUT-X235-LSmitll_NDROT-INt 0 X198-LSmitll_SPLITT-OUT-X235-LSmitll_NDROT-IN 0 z0=5 td=2.6ps
X198 X76-LSmitll_SPLITT-OUT-X198-LSmitll_SPLITT-IN X198-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-INt X198-LSmitll_SPLITT-OUT-X235-LSmitll_NDROT-INt LSmitll_SPLITT

t1173 X199-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt 0 X199-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
t1174 X199-LSmitll_SPLITT-OUT-X237-LSmitll_NDROT-INt 0 X199-LSmitll_SPLITT-OUT-X237-LSmitll_NDROT-IN 0 z0=5 td=1.0ps
X199 X112-LSmitll_SPLITT-OUT-X199-LSmitll_SPLITT-IN X199-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt X199-LSmitll_SPLITT-OUT-X237-LSmitll_NDROT-INt LSmitll_SPLITT

t1175 X200-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt 0 X200-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1176 X200-LSmitll_SPLITT-OUT-X239-LSmitll_NDROT-INt 0 X200-LSmitll_SPLITT-OUT-X239-LSmitll_NDROT-IN 0 z0=5 td=4.1ps
X200 X152-LSmitll_SPLITT-OUT-X200-LSmitll_SPLITT-IN X200-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt X200-LSmitll_SPLITT-OUT-X239-LSmitll_NDROT-INt LSmitll_SPLITT

t1177 X201-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-INt 0 X201-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-IN 0 z0=5 td=4.5ps
t1178 X201-LSmitll_SPLITT-OUT-X241-LSmitll_NDROT-INt 0 X201-LSmitll_SPLITT-OUT-X241-LSmitll_NDROT-IN 0 z0=5 td=1.0ps
X201 X172-LSmitll_SPLITT-OUT-X201-LSmitll_SPLITT-IN X201-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-INt X201-LSmitll_SPLITT-OUT-X241-LSmitll_NDROT-INt LSmitll_SPLITT

t1179 X202-LSmitll_SPLITT-OUT-X244-LSmitll_AND2T-INt 0 X202-LSmitll_SPLITT-OUT-X244-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1180 X202-LSmitll_SPLITT-OUT-X243-LSmitll_NDROT-INt 0 X202-LSmitll_SPLITT-OUT-X243-LSmitll_NDROT-IN 0 z0=5 td=2.3ps
X202 X182-LSmitll_DFFT-OUT-X202-LSmitll_SPLITT-IN X202-LSmitll_SPLITT-OUT-X244-LSmitll_AND2T-INt X202-LSmitll_SPLITT-OUT-X243-LSmitll_NDROT-INt LSmitll_SPLITT

t1181 X203-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-INt 0 X203-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1182 X203-LSmitll_SPLITT-OUT-X245-LSmitll_NDROT-INt 0 X203-LSmitll_SPLITT-OUT-X245-LSmitll_NDROT-IN 0 z0=5 td=1.0ps
X203 X5-LSmitll_SPLITT-OUT-X203-LSmitll_SPLITT-IN X203-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-INt X203-LSmitll_SPLITT-OUT-X245-LSmitll_NDROT-INt LSmitll_SPLITT

t1183 X204-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-INt 0 X204-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1184 X204-LSmitll_SPLITT-OUT-X247-LSmitll_NDROT-INt 0 X204-LSmitll_SPLITT-OUT-X247-LSmitll_NDROT-IN 0 z0=5 td=1.0ps
X204 X46-LSmitll_SPLITT-OUT-X204-LSmitll_SPLITT-IN X204-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-INt X204-LSmitll_SPLITT-OUT-X247-LSmitll_NDROT-INt LSmitll_SPLITT

t1185 X205-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-INt 0 X205-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-IN 0 z0=5 td=3.3ps
t1186 X205-LSmitll_SPLITT-OUT-X249-LSmitll_NDROT-INt 0 X205-LSmitll_SPLITT-OUT-X249-LSmitll_NDROT-IN 0 z0=5 td=1.0ps
X205 X78-LSmitll_SPLITT-OUT-X205-LSmitll_SPLITT-IN X205-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-INt X205-LSmitll_SPLITT-OUT-X249-LSmitll_NDROT-INt LSmitll_SPLITT

t1187 X206-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-INt 0 X206-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-IN 0 z0=5 td=3.2ps
t1188 X206-LSmitll_SPLITT-OUT-X251-LSmitll_NDROT-INt 0 X206-LSmitll_SPLITT-OUT-X251-LSmitll_NDROT-IN 0 z0=5 td=2.3ps
X206 X114-LSmitll_SPLITT-OUT-X206-LSmitll_SPLITT-IN X206-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-INt X206-LSmitll_SPLITT-OUT-X251-LSmitll_NDROT-INt LSmitll_SPLITT

t1189 X207-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-INt 0 X207-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-IN 0 z0=5 td=3.3ps
t1190 X207-LSmitll_SPLITT-OUT-X253-LSmitll_NDROT-INt 0 X207-LSmitll_SPLITT-OUT-X253-LSmitll_NDROT-IN 0 z0=5 td=1.0ps
X207 X154-LSmitll_SPLITT-OUT-X207-LSmitll_SPLITT-IN X207-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-INt X207-LSmitll_SPLITT-OUT-X253-LSmitll_NDROT-INt LSmitll_SPLITT

t1191 X208-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-INt 0 X208-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1192 X208-LSmitll_SPLITT-OUT-X255-LSmitll_NDROT-INt 0 X208-LSmitll_SPLITT-OUT-X255-LSmitll_NDROT-IN 0 z0=5 td=1.0ps
X208 X174-LSmitll_SPLITT-OUT-X208-LSmitll_SPLITT-IN X208-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-INt X208-LSmitll_SPLITT-OUT-X255-LSmitll_NDROT-INt LSmitll_SPLITT

t1193 X209-LSmitll_SPLITT-OUT-X258-LSmitll_AND2T-INt 0 X209-LSmitll_SPLITT-OUT-X258-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t1194 X209-LSmitll_SPLITT-OUT-X257-LSmitll_NDROT-INt 0 X209-LSmitll_SPLITT-OUT-X257-LSmitll_NDROT-IN 0 z0=5 td=2.6ps
X209 X185-LSmitll_DFFT-OUT-X209-LSmitll_SPLITT-IN X209-LSmitll_SPLITT-OUT-X258-LSmitll_AND2T-INt X209-LSmitll_SPLITT-OUT-X257-LSmitll_NDROT-INt LSmitll_SPLITT

t1195 X210-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-INt 0 X210-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t1196 X210-LSmitll_SPLITT-OUT-X259-LSmitll_NDROT-INt 0 X210-LSmitll_SPLITT-OUT-X259-LSmitll_NDROT-IN 0 z0=5 td=2.3ps
X210 X7-LSmitll_SPLITT-OUT-X210-LSmitll_SPLITT-IN X210-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-INt X210-LSmitll_SPLITT-OUT-X259-LSmitll_NDROT-INt LSmitll_SPLITT

t1197 X211-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-INt 0 X211-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
t1198 X211-LSmitll_SPLITT-OUT-X261-LSmitll_NDROT-INt 0 X211-LSmitll_SPLITT-OUT-X261-LSmitll_NDROT-IN 0 z0=5 td=3.6ps
X211 X48-LSmitll_SPLITT-OUT-X211-LSmitll_SPLITT-IN X211-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-INt X211-LSmitll_SPLITT-OUT-X261-LSmitll_NDROT-INt LSmitll_SPLITT

t1199 X212-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-INt 0 X212-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-IN 0 z0=5 td=1.4ps
t1200 X212-LSmitll_SPLITT-OUT-X263-LSmitll_NDROT-INt 0 X212-LSmitll_SPLITT-OUT-X263-LSmitll_NDROT-IN 0 z0=5 td=3.9ps
X212 X80-LSmitll_SPLITT-OUT-X212-LSmitll_SPLITT-IN X212-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-INt X212-LSmitll_SPLITT-OUT-X263-LSmitll_NDROT-INt LSmitll_SPLITT

t1201 X213-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt 0 X213-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
t1202 X213-LSmitll_SPLITT-OUT-X265-LSmitll_NDROT-INt 0 X213-LSmitll_SPLITT-OUT-X265-LSmitll_NDROT-IN 0 z0=5 td=4.1ps
X213 X116-LSmitll_SPLITT-OUT-X213-LSmitll_SPLITT-IN X213-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt X213-LSmitll_SPLITT-OUT-X265-LSmitll_NDROT-INt LSmitll_SPLITT

t1203 X214-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-INt 0 X214-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t1204 X214-LSmitll_SPLITT-OUT-X267-LSmitll_NDROT-INt 0 X214-LSmitll_SPLITT-OUT-X267-LSmitll_NDROT-IN 0 z0=5 td=2.3ps
X214 X156-LSmitll_SPLITT-OUT-X214-LSmitll_SPLITT-IN X214-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-INt X214-LSmitll_SPLITT-OUT-X267-LSmitll_NDROT-INt LSmitll_SPLITT

t1205 X215-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-INt 0 X215-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
t1206 X215-LSmitll_SPLITT-OUT-X269-LSmitll_NDROT-INt 0 X215-LSmitll_SPLITT-OUT-X269-LSmitll_NDROT-IN 0 z0=5 td=2.3ps
X215 X176-LSmitll_SPLITT-OUT-X215-LSmitll_SPLITT-IN X215-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-INt X215-LSmitll_SPLITT-OUT-X269-LSmitll_NDROT-INt LSmitll_SPLITT

t1207 X216-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-INt 0 X216-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-IN 0 z0=5 td=1.4ps
t1208 X216-LSmitll_SPLITT-OUT-X271-LSmitll_NDROT-INt 0 X216-LSmitll_SPLITT-OUT-X271-LSmitll_NDROT-IN 0 z0=5 td=3.1ps
X216 X188-LSmitll_DFFT-OUT-X216-LSmitll_SPLITT-IN X216-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-INt X216-LSmitll_SPLITT-OUT-X271-LSmitll_NDROT-INt LSmitll_SPLITT

t1209 X217-LSmitll_NDROT-OUT-X273-LSmitll_AND2T-INt 0 X217-LSmitll_NDROT-OUT-X273-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X217 X218-LSmitll_AND2T-OUT-X217-LSmitll_NDROT-IN X189-LSmitll_SPLITT-OUT-X217-LSmitll_NDROT-IN X450-LSmitll_SPLITT-OUT-X217-LSmitll_NDROT-IN X217-LSmitll_NDROT-OUT-X273-LSmitll_AND2T-INt LSmitll_NDROT

t1210 X218-LSmitll_AND2T-OUT-X217-LSmitll_NDROT-INt 0 X218-LSmitll_AND2T-OUT-X217-LSmitll_NDROT-IN 0 z0=5 td=3.6ps
X218 X2-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-IN X189-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-IN X455-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-IN X218-LSmitll_AND2T-OUT-X217-LSmitll_NDROT-INt LSmitll_AND2T

t1211 X219-LSmitll_NDROT-OUT-X277-LSmitll_AND2T-INt 0 X219-LSmitll_NDROT-OUT-X277-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
X219 X220-LSmitll_AND2T-OUT-X219-LSmitll_NDROT-IN X190-LSmitll_SPLITT-OUT-X219-LSmitll_NDROT-IN X449-LSmitll_SPLITT-OUT-X219-LSmitll_NDROT-IN X219-LSmitll_NDROT-OUT-X277-LSmitll_AND2T-INt LSmitll_NDROT

t1212 X220-LSmitll_AND2T-OUT-X219-LSmitll_NDROT-INt 0 X220-LSmitll_AND2T-OUT-X219-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
X220 X41-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-IN X190-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-IN X547-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-IN X220-LSmitll_AND2T-OUT-X219-LSmitll_NDROT-INt LSmitll_AND2T

t1213 X221-LSmitll_NDROT-OUT-X281-LSmitll_AND2T-INt 0 X221-LSmitll_NDROT-OUT-X281-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X221 X222-LSmitll_AND2T-OUT-X221-LSmitll_NDROT-IN X191-LSmitll_SPLITT-OUT-X221-LSmitll_NDROT-IN X548-LSmitll_SPLITT-OUT-X221-LSmitll_NDROT-IN X221-LSmitll_NDROT-OUT-X281-LSmitll_AND2T-INt LSmitll_NDROT

t1214 X222-LSmitll_AND2T-OUT-X221-LSmitll_NDROT-INt 0 X222-LSmitll_AND2T-OUT-X221-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
X222 X73-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-IN X191-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-IN X466-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-IN X222-LSmitll_AND2T-OUT-X221-LSmitll_NDROT-INt LSmitll_AND2T

t1215 X223-LSmitll_NDROT-OUT-X285-LSmitll_AND2T-INt 0 X223-LSmitll_NDROT-OUT-X285-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X223 X224-LSmitll_AND2T-OUT-X223-LSmitll_NDROT-IN X192-LSmitll_SPLITT-OUT-X223-LSmitll_NDROT-IN X549-LSmitll_SPLITT-OUT-X223-LSmitll_NDROT-IN X223-LSmitll_NDROT-OUT-X285-LSmitll_AND2T-INt LSmitll_NDROT

t1216 X224-LSmitll_AND2T-OUT-X223-LSmitll_NDROT-INt 0 X224-LSmitll_AND2T-OUT-X223-LSmitll_NDROT-IN 0 z0=5 td=2.4ps
X224 X109-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-IN X192-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-IN X463-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-IN X224-LSmitll_AND2T-OUT-X223-LSmitll_NDROT-INt LSmitll_AND2T

t1217 X225-LSmitll_NDROT-OUT-X289-LSmitll_AND2T-INt 0 X225-LSmitll_NDROT-OUT-X289-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
X225 X226-LSmitll_AND2T-OUT-X225-LSmitll_NDROT-IN X193-LSmitll_SPLITT-OUT-X225-LSmitll_NDROT-IN X499-LSmitll_SPLITT-OUT-X225-LSmitll_NDROT-IN X225-LSmitll_NDROT-OUT-X289-LSmitll_AND2T-INt LSmitll_NDROT

t1218 X226-LSmitll_AND2T-OUT-X225-LSmitll_NDROT-INt 0 X226-LSmitll_AND2T-OUT-X225-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
X226 X149-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-IN X193-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-IN X500-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-IN X226-LSmitll_AND2T-OUT-X225-LSmitll_NDROT-INt LSmitll_AND2T

t1219 X227-LSmitll_NDROT-OUT-X293-LSmitll_AND2T-INt 0 X227-LSmitll_NDROT-OUT-X293-LSmitll_AND2T-IN 0 z0=5 td=2.3ps
X227 X228-LSmitll_AND2T-OUT-X227-LSmitll_NDROT-IN X194-LSmitll_SPLITT-OUT-X227-LSmitll_NDROT-IN X516-LSmitll_SPLITT-OUT-X227-LSmitll_NDROT-IN X227-LSmitll_NDROT-OUT-X293-LSmitll_AND2T-INt LSmitll_NDROT

t1220 X228-LSmitll_AND2T-OUT-X227-LSmitll_NDROT-INt 0 X228-LSmitll_AND2T-OUT-X227-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
X228 X169-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-IN X194-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-IN X550-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-IN X228-LSmitll_AND2T-OUT-X227-LSmitll_NDROT-INt LSmitll_AND2T

t1221 X229-LSmitll_NDROT-OUT-X297-LSmitll_AND2T-INt 0 X229-LSmitll_NDROT-OUT-X297-LSmitll_AND2T-IN 0 z0=5 td=4.8ps
X229 X230-LSmitll_AND2T-OUT-X229-LSmitll_NDROT-IN X195-LSmitll_SPLITT-OUT-X229-LSmitll_NDROT-IN X487-LSmitll_SPLITT-OUT-X229-LSmitll_NDROT-IN X229-LSmitll_NDROT-OUT-X297-LSmitll_AND2T-INt LSmitll_NDROT

t1222 X230-LSmitll_AND2T-OUT-X229-LSmitll_NDROT-INt 0 X230-LSmitll_AND2T-OUT-X229-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
X230 X177-LSmitll_DFFT-OUT-X230-LSmitll_AND2T-IN X195-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-IN X487-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-IN X230-LSmitll_AND2T-OUT-X229-LSmitll_NDROT-INt LSmitll_AND2T

t1223 X231-LSmitll_NDROT-OUT-X274-LSmitll_AND2T-INt 0 X231-LSmitll_NDROT-OUT-X274-LSmitll_AND2T-IN 0 z0=5 td=3.8ps
X231 X232-LSmitll_AND2T-OUT-X231-LSmitll_NDROT-IN X196-LSmitll_SPLITT-OUT-X231-LSmitll_NDROT-IN X425-LSmitll_SPLITT-OUT-X231-LSmitll_NDROT-IN X231-LSmitll_NDROT-OUT-X274-LSmitll_AND2T-INt LSmitll_NDROT

t1224 X232-LSmitll_AND2T-OUT-X231-LSmitll_NDROT-INt 0 X232-LSmitll_AND2T-OUT-X231-LSmitll_NDROT-IN 0 z0=5 td=3.8ps
X232 X4-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-IN X196-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-IN X551-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-IN X232-LSmitll_AND2T-OUT-X231-LSmitll_NDROT-INt LSmitll_AND2T

t1225 X233-LSmitll_NDROT-OUT-X278-LSmitll_AND2T-INt 0 X233-LSmitll_NDROT-OUT-X278-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X233 X234-LSmitll_AND2T-OUT-X233-LSmitll_NDROT-IN X197-LSmitll_SPLITT-OUT-X233-LSmitll_NDROT-IN X355-LSmitll_SPLITT-OUT-X233-LSmitll_NDROT-IN X233-LSmitll_NDROT-OUT-X278-LSmitll_AND2T-INt LSmitll_NDROT

t1226 X234-LSmitll_AND2T-OUT-X233-LSmitll_NDROT-INt 0 X234-LSmitll_AND2T-OUT-X233-LSmitll_NDROT-IN 0 z0=5 td=3.5ps
X234 X43-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN X197-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN X552-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN X234-LSmitll_AND2T-OUT-X233-LSmitll_NDROT-INt LSmitll_AND2T

t1227 X235-LSmitll_NDROT-OUT-X282-LSmitll_AND2T-INt 0 X235-LSmitll_NDROT-OUT-X282-LSmitll_AND2T-IN 0 z0=5 td=3.1ps
X235 X236-LSmitll_AND2T-OUT-X235-LSmitll_NDROT-IN X198-LSmitll_SPLITT-OUT-X235-LSmitll_NDROT-IN X553-LSmitll_SPLITT-OUT-X235-LSmitll_NDROT-IN X235-LSmitll_NDROT-OUT-X282-LSmitll_AND2T-INt LSmitll_NDROT

t1228 X236-LSmitll_AND2T-OUT-X235-LSmitll_NDROT-INt 0 X236-LSmitll_AND2T-OUT-X235-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
X236 X75-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-IN X198-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-IN X444-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-IN X236-LSmitll_AND2T-OUT-X235-LSmitll_NDROT-INt LSmitll_AND2T

t1229 X237-LSmitll_NDROT-OUT-X286-LSmitll_AND2T-INt 0 X237-LSmitll_NDROT-OUT-X286-LSmitll_AND2T-IN 0 z0=5 td=7.4ps
X237 X238-LSmitll_AND2T-OUT-X237-LSmitll_NDROT-IN X199-LSmitll_SPLITT-OUT-X237-LSmitll_NDROT-IN X463-LSmitll_SPLITT-OUT-X237-LSmitll_NDROT-IN X237-LSmitll_NDROT-OUT-X286-LSmitll_AND2T-INt LSmitll_NDROT

t1230 X238-LSmitll_AND2T-OUT-X237-LSmitll_NDROT-INt 0 X238-LSmitll_AND2T-OUT-X237-LSmitll_NDROT-IN 0 z0=5 td=2.9ps
X238 X111-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN X199-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN X554-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN X238-LSmitll_AND2T-OUT-X237-LSmitll_NDROT-INt LSmitll_AND2T

t1231 X239-LSmitll_NDROT-OUT-X290-LSmitll_AND2T-INt 0 X239-LSmitll_NDROT-OUT-X290-LSmitll_AND2T-IN 0 z0=5 td=3.1ps
X239 X240-LSmitll_AND2T-OUT-X239-LSmitll_NDROT-IN X200-LSmitll_SPLITT-OUT-X239-LSmitll_NDROT-IN X391-LSmitll_SPLITT-OUT-X239-LSmitll_NDROT-IN X239-LSmitll_NDROT-OUT-X290-LSmitll_AND2T-INt LSmitll_NDROT

t1232 X240-LSmitll_AND2T-OUT-X239-LSmitll_NDROT-INt 0 X240-LSmitll_AND2T-OUT-X239-LSmitll_NDROT-IN 0 z0=5 td=2.9ps
X240 X151-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN X200-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN X386-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN X240-LSmitll_AND2T-OUT-X239-LSmitll_NDROT-INt LSmitll_AND2T

t1233 X241-LSmitll_NDROT-OUT-X294-LSmitll_AND2T-INt 0 X241-LSmitll_NDROT-OUT-X294-LSmitll_AND2T-IN 0 z0=5 td=9.1ps
X241 X242-LSmitll_AND2T-OUT-X241-LSmitll_NDROT-IN X201-LSmitll_SPLITT-OUT-X241-LSmitll_NDROT-IN X518-LSmitll_SPLITT-OUT-X241-LSmitll_NDROT-IN X241-LSmitll_NDROT-OUT-X294-LSmitll_AND2T-INt LSmitll_NDROT

t1234 X242-LSmitll_AND2T-OUT-X241-LSmitll_NDROT-INt 0 X242-LSmitll_AND2T-OUT-X241-LSmitll_NDROT-IN 0 z0=5 td=3.1ps
X242 X171-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-IN X201-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-IN X516-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-IN X242-LSmitll_AND2T-OUT-X241-LSmitll_NDROT-INt LSmitll_AND2T

t1235 X243-LSmitll_NDROT-OUT-X298-LSmitll_AND2T-INt 0 X243-LSmitll_NDROT-OUT-X298-LSmitll_AND2T-IN 0 z0=5 td=3.3ps
X243 X244-LSmitll_AND2T-OUT-X243-LSmitll_NDROT-IN X202-LSmitll_SPLITT-OUT-X243-LSmitll_NDROT-IN X555-LSmitll_SPLITT-OUT-X243-LSmitll_NDROT-IN X243-LSmitll_NDROT-OUT-X298-LSmitll_AND2T-INt LSmitll_NDROT

t1236 X244-LSmitll_AND2T-OUT-X243-LSmitll_NDROT-INt 0 X244-LSmitll_AND2T-OUT-X243-LSmitll_NDROT-IN 0 z0=5 td=2.9ps
X244 X180-LSmitll_DFFT-OUT-X244-LSmitll_AND2T-IN X202-LSmitll_SPLITT-OUT-X244-LSmitll_AND2T-IN X494-LSmitll_SPLITT-OUT-X244-LSmitll_AND2T-IN X244-LSmitll_AND2T-OUT-X243-LSmitll_NDROT-INt LSmitll_AND2T

t1237 X245-LSmitll_NDROT-OUT-X275-LSmitll_AND2T-INt 0 X245-LSmitll_NDROT-OUT-X275-LSmitll_AND2T-IN 0 z0=5 td=3.6ps
X245 X246-LSmitll_AND2T-OUT-X245-LSmitll_NDROT-IN X203-LSmitll_SPLITT-OUT-X245-LSmitll_NDROT-IN X556-LSmitll_SPLITT-OUT-X245-LSmitll_NDROT-IN X245-LSmitll_NDROT-OUT-X275-LSmitll_AND2T-INt LSmitll_NDROT

t1238 X246-LSmitll_AND2T-OUT-X245-LSmitll_NDROT-INt 0 X246-LSmitll_AND2T-OUT-X245-LSmitll_NDROT-IN 0 z0=5 td=2.4ps
X246 X6-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-IN X203-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-IN X424-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-IN X246-LSmitll_AND2T-OUT-X245-LSmitll_NDROT-INt LSmitll_AND2T

t1239 X247-LSmitll_NDROT-OUT-X279-LSmitll_AND2T-INt 0 X247-LSmitll_NDROT-OUT-X279-LSmitll_AND2T-IN 0 z0=5 td=5.1ps
X247 X248-LSmitll_AND2T-OUT-X247-LSmitll_NDROT-IN X204-LSmitll_SPLITT-OUT-X247-LSmitll_NDROT-IN X330-LSmitll_SPLITT-OUT-X247-LSmitll_NDROT-IN X247-LSmitll_NDROT-OUT-X279-LSmitll_AND2T-INt LSmitll_NDROT

t1240 X248-LSmitll_AND2T-OUT-X247-LSmitll_NDROT-INt 0 X248-LSmitll_AND2T-OUT-X247-LSmitll_NDROT-IN 0 z0=5 td=2.4ps
X248 X45-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-IN X204-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-IN X347-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-IN X248-LSmitll_AND2T-OUT-X247-LSmitll_NDROT-INt LSmitll_AND2T

t1241 X249-LSmitll_NDROT-OUT-X283-LSmitll_AND2T-INt 0 X249-LSmitll_NDROT-OUT-X283-LSmitll_AND2T-IN 0 z0=5 td=3.6ps
X249 X250-LSmitll_AND2T-OUT-X249-LSmitll_NDROT-IN X205-LSmitll_SPLITT-OUT-X249-LSmitll_NDROT-IN X360-LSmitll_SPLITT-OUT-X249-LSmitll_NDROT-IN X249-LSmitll_NDROT-OUT-X283-LSmitll_AND2T-INt LSmitll_NDROT

t1242 X250-LSmitll_AND2T-OUT-X249-LSmitll_NDROT-INt 0 X250-LSmitll_AND2T-OUT-X249-LSmitll_NDROT-IN 0 z0=5 td=12.3ps
X250 X77-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-IN X205-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-IN X557-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-IN X250-LSmitll_AND2T-OUT-X249-LSmitll_NDROT-INt LSmitll_AND2T

t1243 X251-LSmitll_NDROT-OUT-X287-LSmitll_AND2T-INt 0 X251-LSmitll_NDROT-OUT-X287-LSmitll_AND2T-IN 0 z0=5 td=4.9ps
X251 X252-LSmitll_AND2T-OUT-X251-LSmitll_NDROT-IN X206-LSmitll_SPLITT-OUT-X251-LSmitll_NDROT-IN X367-LSmitll_SPLITT-OUT-X251-LSmitll_NDROT-IN X251-LSmitll_NDROT-OUT-X287-LSmitll_AND2T-INt LSmitll_NDROT

t1244 X252-LSmitll_AND2T-OUT-X251-LSmitll_NDROT-INt 0 X252-LSmitll_AND2T-OUT-X251-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
X252 X113-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-IN X206-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-IN X558-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-IN X252-LSmitll_AND2T-OUT-X251-LSmitll_NDROT-INt LSmitll_AND2T

t1245 X253-LSmitll_NDROT-OUT-X291-LSmitll_AND2T-INt 0 X253-LSmitll_NDROT-OUT-X291-LSmitll_AND2T-IN 0 z0=5 td=1.1ps
X253 X254-LSmitll_AND2T-OUT-X253-LSmitll_NDROT-IN X207-LSmitll_SPLITT-OUT-X253-LSmitll_NDROT-IN X559-LSmitll_SPLITT-OUT-X253-LSmitll_NDROT-IN X253-LSmitll_NDROT-OUT-X291-LSmitll_AND2T-INt LSmitll_NDROT

t1246 X254-LSmitll_AND2T-OUT-X253-LSmitll_NDROT-INt 0 X254-LSmitll_AND2T-OUT-X253-LSmitll_NDROT-IN 0 z0=5 td=3.5ps
X254 X153-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-IN X207-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-IN X474-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-IN X254-LSmitll_AND2T-OUT-X253-LSmitll_NDROT-INt LSmitll_AND2T

t1247 X255-LSmitll_NDROT-OUT-X295-LSmitll_AND2T-INt 0 X255-LSmitll_NDROT-OUT-X295-LSmitll_AND2T-IN 0 z0=5 td=4.1ps
X255 X256-LSmitll_AND2T-OUT-X255-LSmitll_NDROT-IN X208-LSmitll_SPLITT-OUT-X255-LSmitll_NDROT-IN X477-LSmitll_SPLITT-OUT-X255-LSmitll_NDROT-IN X255-LSmitll_NDROT-OUT-X295-LSmitll_AND2T-INt LSmitll_NDROT

t1248 X256-LSmitll_AND2T-OUT-X255-LSmitll_NDROT-INt 0 X256-LSmitll_AND2T-OUT-X255-LSmitll_NDROT-IN 0 z0=5 td=2.4ps
X256 X173-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-IN X208-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-IN X477-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-IN X256-LSmitll_AND2T-OUT-X255-LSmitll_NDROT-INt LSmitll_AND2T

t1249 X257-LSmitll_NDROT-OUT-X299-LSmitll_AND2T-INt 0 X257-LSmitll_NDROT-OUT-X299-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X257 X258-LSmitll_AND2T-OUT-X257-LSmitll_NDROT-IN X209-LSmitll_SPLITT-OUT-X257-LSmitll_NDROT-IN X560-LSmitll_SPLITT-OUT-X257-LSmitll_NDROT-IN X257-LSmitll_NDROT-OUT-X299-LSmitll_AND2T-INt LSmitll_NDROT

t1250 X258-LSmitll_AND2T-OUT-X257-LSmitll_NDROT-INt 0 X258-LSmitll_AND2T-OUT-X257-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
X258 X183-LSmitll_DFFT-OUT-X258-LSmitll_AND2T-IN X209-LSmitll_SPLITT-OUT-X258-LSmitll_AND2T-IN X561-LSmitll_SPLITT-OUT-X258-LSmitll_AND2T-IN X258-LSmitll_AND2T-OUT-X257-LSmitll_NDROT-INt LSmitll_AND2T

t1251 X259-LSmitll_NDROT-OUT-X276-LSmitll_AND2T-INt 0 X259-LSmitll_NDROT-OUT-X276-LSmitll_AND2T-IN 0 z0=5 td=11.2ps
X259 X260-LSmitll_AND2T-OUT-X259-LSmitll_NDROT-IN X210-LSmitll_SPLITT-OUT-X259-LSmitll_NDROT-IN X347-LSmitll_SPLITT-OUT-X259-LSmitll_NDROT-IN X259-LSmitll_NDROT-OUT-X276-LSmitll_AND2T-INt LSmitll_NDROT

t1252 X260-LSmitll_AND2T-OUT-X259-LSmitll_NDROT-INt 0 X260-LSmitll_AND2T-OUT-X259-LSmitll_NDROT-IN 0 z0=5 td=4.2ps
X260 X8-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-IN X210-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-IN X562-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-IN X260-LSmitll_AND2T-OUT-X259-LSmitll_NDROT-INt LSmitll_AND2T

t1253 X261-LSmitll_NDROT-OUT-X280-LSmitll_AND2T-INt 0 X261-LSmitll_NDROT-OUT-X280-LSmitll_AND2T-IN 0 z0=5 td=4.0ps
X261 X262-LSmitll_AND2T-OUT-X261-LSmitll_NDROT-IN X211-LSmitll_SPLITT-OUT-X261-LSmitll_NDROT-IN X322-LSmitll_SPLITT-OUT-X261-LSmitll_NDROT-IN X261-LSmitll_NDROT-OUT-X280-LSmitll_AND2T-INt LSmitll_NDROT

t1254 X262-LSmitll_AND2T-OUT-X261-LSmitll_NDROT-INt 0 X262-LSmitll_AND2T-OUT-X261-LSmitll_NDROT-IN 0 z0=5 td=2.9ps
X262 X47-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-IN X211-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-IN X322-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-IN X262-LSmitll_AND2T-OUT-X261-LSmitll_NDROT-INt LSmitll_AND2T

t1255 X263-LSmitll_NDROT-OUT-X284-LSmitll_AND2T-INt 0 X263-LSmitll_NDROT-OUT-X284-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
X263 X264-LSmitll_AND2T-OUT-X263-LSmitll_NDROT-IN X212-LSmitll_SPLITT-OUT-X263-LSmitll_NDROT-IN X563-LSmitll_SPLITT-OUT-X263-LSmitll_NDROT-IN X263-LSmitll_NDROT-OUT-X284-LSmitll_AND2T-INt LSmitll_NDROT

t1256 X264-LSmitll_AND2T-OUT-X263-LSmitll_NDROT-INt 0 X264-LSmitll_AND2T-OUT-X263-LSmitll_NDROT-IN 0 z0=5 td=2.9ps
X264 X79-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-IN X212-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-IN X340-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-IN X264-LSmitll_AND2T-OUT-X263-LSmitll_NDROT-INt LSmitll_AND2T

t1257 X265-LSmitll_NDROT-OUT-X288-LSmitll_AND2T-INt 0 X265-LSmitll_NDROT-OUT-X288-LSmitll_AND2T-IN 0 z0=5 td=2.7ps
X265 X266-LSmitll_AND2T-OUT-X265-LSmitll_NDROT-IN X213-LSmitll_SPLITT-OUT-X265-LSmitll_NDROT-IN X342-LSmitll_SPLITT-OUT-X265-LSmitll_NDROT-IN X265-LSmitll_NDROT-OUT-X288-LSmitll_AND2T-INt LSmitll_NDROT

t1258 X266-LSmitll_AND2T-OUT-X265-LSmitll_NDROT-INt 0 X266-LSmitll_AND2T-OUT-X265-LSmitll_NDROT-IN 0 z0=5 td=3.3ps
X266 X115-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN X213-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN X342-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN X266-LSmitll_AND2T-OUT-X265-LSmitll_NDROT-INt LSmitll_AND2T

t1259 X267-LSmitll_NDROT-OUT-X292-LSmitll_AND2T-INt 0 X267-LSmitll_NDROT-OUT-X292-LSmitll_AND2T-IN 0 z0=5 td=2.7ps
X267 X268-LSmitll_AND2T-OUT-X267-LSmitll_NDROT-IN X214-LSmitll_SPLITT-OUT-X267-LSmitll_NDROT-IN X399-LSmitll_SPLITT-OUT-X267-LSmitll_NDROT-IN X267-LSmitll_NDROT-OUT-X292-LSmitll_AND2T-INt LSmitll_NDROT

t1260 X268-LSmitll_AND2T-OUT-X267-LSmitll_NDROT-INt 0 X268-LSmitll_AND2T-OUT-X267-LSmitll_NDROT-IN 0 z0=5 td=4.0ps
X268 X155-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-IN X214-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-IN X398-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-IN X268-LSmitll_AND2T-OUT-X267-LSmitll_NDROT-INt LSmitll_AND2T

t1261 X269-LSmitll_NDROT-OUT-X296-LSmitll_AND2T-INt 0 X269-LSmitll_NDROT-OUT-X296-LSmitll_AND2T-IN 0 z0=5 td=2.6ps
X269 X270-LSmitll_AND2T-OUT-X269-LSmitll_NDROT-IN X215-LSmitll_SPLITT-OUT-X269-LSmitll_NDROT-IN X401-LSmitll_SPLITT-OUT-X269-LSmitll_NDROT-IN X269-LSmitll_NDROT-OUT-X296-LSmitll_AND2T-INt LSmitll_NDROT

t1262 X270-LSmitll_AND2T-OUT-X269-LSmitll_NDROT-INt 0 X270-LSmitll_AND2T-OUT-X269-LSmitll_NDROT-IN 0 z0=5 td=5.4ps
X270 X175-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-IN X215-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-IN X381-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-IN X270-LSmitll_AND2T-OUT-X269-LSmitll_NDROT-INt LSmitll_AND2T

t1263 X271-LSmitll_NDROT-OUT-X300-LSmitll_AND2T-INt 0 X271-LSmitll_NDROT-OUT-X300-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
X271 X272-LSmitll_AND2T-OUT-X271-LSmitll_NDROT-IN X216-LSmitll_SPLITT-OUT-X271-LSmitll_NDROT-IN X564-LSmitll_SPLITT-OUT-X271-LSmitll_NDROT-IN X271-LSmitll_NDROT-OUT-X300-LSmitll_AND2T-INt LSmitll_NDROT

t1264 X272-LSmitll_AND2T-OUT-X271-LSmitll_NDROT-INt 0 X272-LSmitll_AND2T-OUT-X271-LSmitll_NDROT-IN 0 z0=5 td=3.1ps
X272 X186-LSmitll_DFFT-OUT-X272-LSmitll_AND2T-IN X216-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-IN X386-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-IN X272-LSmitll_AND2T-OUT-X271-LSmitll_NDROT-INt LSmitll_AND2T

t1265 X273-LSmitll_AND2T-OUT-X301-LSmitll_OR2T-INt 0 X273-LSmitll_AND2T-OUT-X301-LSmitll_OR2T-IN 0 z0=5 td=12.7ps
X273 X217-LSmitll_NDROT-OUT-X273-LSmitll_AND2T-IN X130-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-IN X449-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-IN X273-LSmitll_AND2T-OUT-X301-LSmitll_OR2T-INt LSmitll_AND2T

t1266 X274-LSmitll_AND2T-OUT-X301-LSmitll_OR2T-INt 0 X274-LSmitll_AND2T-OUT-X301-LSmitll_OR2T-IN 0 z0=5 td=1.3ps
X274 X231-LSmitll_NDROT-OUT-X274-LSmitll_AND2T-IN X128-LSmitll_SPLITT-OUT-X274-LSmitll_AND2T-IN X424-LSmitll_SPLITT-OUT-X274-LSmitll_AND2T-IN X274-LSmitll_AND2T-OUT-X301-LSmitll_OR2T-INt LSmitll_AND2T

t1267 X275-LSmitll_AND2T-OUT-X302-LSmitll_OR2T-INt 0 X275-LSmitll_AND2T-OUT-X302-LSmitll_OR2T-IN 0 z0=5 td=0.9ps
X275 X245-LSmitll_NDROT-OUT-X275-LSmitll_AND2T-IN X127-LSmitll_SPLITT-OUT-X275-LSmitll_AND2T-IN X353-LSmitll_SPLITT-OUT-X275-LSmitll_AND2T-IN X275-LSmitll_AND2T-OUT-X302-LSmitll_OR2T-INt LSmitll_AND2T

t1268 X276-LSmitll_AND2T-OUT-X302-LSmitll_OR2T-INt 0 X276-LSmitll_AND2T-OUT-X302-LSmitll_OR2T-IN 0 z0=5 td=14.7ps
X276 X259-LSmitll_NDROT-OUT-X276-LSmitll_AND2T-IN X125-LSmitll_SPLITT-OUT-X276-LSmitll_AND2T-IN X328-LSmitll_SPLITT-OUT-X276-LSmitll_AND2T-IN X276-LSmitll_AND2T-OUT-X302-LSmitll_OR2T-INt LSmitll_AND2T

t1269 X277-LSmitll_AND2T-OUT-X303-LSmitll_OR2T-INt 0 X277-LSmitll_AND2T-OUT-X303-LSmitll_OR2T-IN 0 z0=5 td=4.6ps
X277 X130-LSmitll_SPLITT-OUT-X277-LSmitll_AND2T-IN X219-LSmitll_NDROT-OUT-X277-LSmitll_AND2T-IN X565-LSmitll_SPLITT-OUT-X277-LSmitll_AND2T-IN X277-LSmitll_AND2T-OUT-X303-LSmitll_OR2T-INt LSmitll_AND2T

t1270 X278-LSmitll_AND2T-OUT-X303-LSmitll_OR2T-INt 0 X278-LSmitll_AND2T-OUT-X303-LSmitll_OR2T-IN 0 z0=5 td=19.1ps
X278 X128-LSmitll_SPLITT-OUT-X278-LSmitll_AND2T-IN X233-LSmitll_NDROT-OUT-X278-LSmitll_AND2T-IN X355-LSmitll_SPLITT-OUT-X278-LSmitll_AND2T-IN X278-LSmitll_AND2T-OUT-X303-LSmitll_OR2T-INt LSmitll_AND2T

t1271 X279-LSmitll_AND2T-OUT-X304-LSmitll_OR2T-INt 0 X279-LSmitll_AND2T-OUT-X304-LSmitll_OR2T-IN 0 z0=5 td=2.4ps
X279 X127-LSmitll_SPLITT-OUT-X279-LSmitll_AND2T-IN X247-LSmitll_NDROT-OUT-X279-LSmitll_AND2T-IN X350-LSmitll_SPLITT-OUT-X279-LSmitll_AND2T-IN X279-LSmitll_AND2T-OUT-X304-LSmitll_OR2T-INt LSmitll_AND2T

t1272 X280-LSmitll_AND2T-OUT-X304-LSmitll_OR2T-INt 0 X280-LSmitll_AND2T-OUT-X304-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X280 X125-LSmitll_SPLITT-OUT-X280-LSmitll_AND2T-IN X261-LSmitll_NDROT-OUT-X280-LSmitll_AND2T-IN X566-LSmitll_SPLITT-OUT-X280-LSmitll_AND2T-IN X280-LSmitll_AND2T-OUT-X304-LSmitll_OR2T-INt LSmitll_AND2T

t1273 X281-LSmitll_AND2T-OUT-X305-LSmitll_OR2T-INt 0 X281-LSmitll_AND2T-OUT-X305-LSmitll_OR2T-IN 0 z0=5 td=12.0ps
X281 X120-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-IN X221-LSmitll_NDROT-OUT-X281-LSmitll_AND2T-IN X461-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-IN X281-LSmitll_AND2T-OUT-X305-LSmitll_OR2T-INt LSmitll_AND2T

t1274 X282-LSmitll_AND2T-OUT-X305-LSmitll_OR2T-INt 0 X282-LSmitll_AND2T-OUT-X305-LSmitll_OR2T-IN 0 z0=5 td=1.3ps
X282 X235-LSmitll_NDROT-OUT-X282-LSmitll_AND2T-IN X129-LSmitll_SPLITT-OUT-X282-LSmitll_AND2T-IN X437-LSmitll_SPLITT-OUT-X282-LSmitll_AND2T-IN X282-LSmitll_AND2T-OUT-X305-LSmitll_OR2T-INt LSmitll_AND2T

t1275 X283-LSmitll_AND2T-OUT-X306-LSmitll_OR2T-INt 0 X283-LSmitll_AND2T-OUT-X306-LSmitll_OR2T-IN 0 z0=5 td=20.2ps
X283 X118-LSmitll_SPLITT-OUT-X283-LSmitll_AND2T-IN X249-LSmitll_NDROT-OUT-X283-LSmitll_AND2T-IN X567-LSmitll_SPLITT-OUT-X283-LSmitll_AND2T-IN X283-LSmitll_AND2T-OUT-X306-LSmitll_OR2T-INt LSmitll_AND2T

t1276 X284-LSmitll_AND2T-OUT-X306-LSmitll_OR2T-INt 0 X284-LSmitll_AND2T-OUT-X306-LSmitll_OR2T-IN 0 z0=5 td=4.0ps
X284 X263-LSmitll_NDROT-OUT-X284-LSmitll_AND2T-IN X126-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-IN X340-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-IN X284-LSmitll_AND2T-OUT-X306-LSmitll_OR2T-INt LSmitll_AND2T

t1277 X285-LSmitll_AND2T-OUT-X307-LSmitll_OR2T-INt 0 X285-LSmitll_AND2T-OUT-X307-LSmitll_OR2T-IN 0 z0=5 td=0.9ps
X285 X223-LSmitll_NDROT-OUT-X285-LSmitll_AND2T-IN X135-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-IN X480-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-IN X285-LSmitll_AND2T-OUT-X307-LSmitll_OR2T-INt LSmitll_AND2T

t1278 X286-LSmitll_AND2T-OUT-X307-LSmitll_OR2T-INt 0 X286-LSmitll_AND2T-OUT-X307-LSmitll_OR2T-IN 0 z0=5 td=2.3ps
X286 X129-LSmitll_SPLITT-OUT-X286-LSmitll_AND2T-IN X237-LSmitll_NDROT-OUT-X286-LSmitll_AND2T-IN X444-LSmitll_SPLITT-OUT-X286-LSmitll_AND2T-IN X286-LSmitll_AND2T-OUT-X307-LSmitll_OR2T-INt LSmitll_AND2T

t1279 X287-LSmitll_AND2T-OUT-X308-LSmitll_OR2T-INt 0 X287-LSmitll_AND2T-OUT-X308-LSmitll_OR2T-IN 0 z0=5 td=8.7ps
X287 X251-LSmitll_NDROT-OUT-X287-LSmitll_AND2T-IN X132-LSmitll_SPLITT-OUT-X287-LSmitll_AND2T-IN X404-LSmitll_SPLITT-OUT-X287-LSmitll_AND2T-IN X287-LSmitll_AND2T-OUT-X308-LSmitll_OR2T-INt LSmitll_AND2T

t1280 X288-LSmitll_AND2T-OUT-X308-LSmitll_OR2T-INt 0 X288-LSmitll_AND2T-OUT-X308-LSmitll_OR2T-IN 0 z0=5 td=12.0ps
X288 X126-LSmitll_SPLITT-OUT-X288-LSmitll_AND2T-IN X265-LSmitll_NDROT-OUT-X288-LSmitll_AND2T-IN X362-LSmitll_SPLITT-OUT-X288-LSmitll_AND2T-IN X288-LSmitll_AND2T-OUT-X308-LSmitll_OR2T-INt LSmitll_AND2T

t1281 X289-LSmitll_AND2T-OUT-X309-LSmitll_OR2T-INt 0 X289-LSmitll_AND2T-OUT-X309-LSmitll_OR2T-IN 0 z0=5 td=16.1ps
X289 X135-LSmitll_SPLITT-OUT-X289-LSmitll_AND2T-IN X225-LSmitll_NDROT-OUT-X289-LSmitll_AND2T-IN X499-LSmitll_SPLITT-OUT-X289-LSmitll_AND2T-IN X289-LSmitll_AND2T-OUT-X309-LSmitll_OR2T-INt LSmitll_AND2T

t1282 X290-LSmitll_AND2T-OUT-X309-LSmitll_OR2T-INt 0 X290-LSmitll_AND2T-OUT-X309-LSmitll_OR2T-IN 0 z0=5 td=17.7ps
X290 X239-LSmitll_NDROT-OUT-X290-LSmitll_AND2T-IN X134-LSmitll_SPLITT-OUT-X290-LSmitll_AND2T-IN X391-LSmitll_SPLITT-OUT-X290-LSmitll_AND2T-IN X290-LSmitll_AND2T-OUT-X309-LSmitll_OR2T-INt LSmitll_AND2T

t1283 X291-LSmitll_AND2T-OUT-X310-LSmitll_OR2T-INt 0 X291-LSmitll_AND2T-OUT-X310-LSmitll_OR2T-IN 0 z0=5 td=0.9ps
X291 X132-LSmitll_SPLITT-OUT-X291-LSmitll_AND2T-IN X253-LSmitll_NDROT-OUT-X291-LSmitll_AND2T-IN X406-LSmitll_SPLITT-OUT-X291-LSmitll_AND2T-IN X291-LSmitll_AND2T-OUT-X310-LSmitll_OR2T-INt LSmitll_AND2T

t1284 X292-LSmitll_AND2T-OUT-X310-LSmitll_OR2T-INt 0 X292-LSmitll_AND2T-OUT-X310-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X292 X267-LSmitll_NDROT-OUT-X292-LSmitll_AND2T-IN X131-LSmitll_SPLITT-OUT-X292-LSmitll_AND2T-IN X401-LSmitll_SPLITT-OUT-X292-LSmitll_AND2T-IN X292-LSmitll_AND2T-OUT-X310-LSmitll_OR2T-INt LSmitll_AND2T

t1285 X293-LSmitll_AND2T-OUT-X311-LSmitll_OR2T-INt 0 X293-LSmitll_AND2T-OUT-X311-LSmitll_OR2T-IN 0 z0=5 td=2.5ps
X293 X227-LSmitll_NDROT-OUT-X293-LSmitll_AND2T-IN X136-LSmitll_SPLITT-OUT-X293-LSmitll_AND2T-IN X415-LSmitll_SPLITT-OUT-X293-LSmitll_AND2T-IN X293-LSmitll_AND2T-OUT-X311-LSmitll_OR2T-INt LSmitll_AND2T

t1286 X294-LSmitll_AND2T-OUT-X311-LSmitll_OR2T-INt 0 X294-LSmitll_AND2T-OUT-X311-LSmitll_OR2T-IN 0 z0=5 td=10.2ps
X294 X134-LSmitll_SPLITT-OUT-X294-LSmitll_AND2T-IN X241-LSmitll_NDROT-OUT-X294-LSmitll_AND2T-IN X492-LSmitll_SPLITT-OUT-X294-LSmitll_AND2T-IN X294-LSmitll_AND2T-OUT-X311-LSmitll_OR2T-INt LSmitll_AND2T

t1287 X295-LSmitll_AND2T-OUT-X312-LSmitll_OR2T-INt 0 X295-LSmitll_AND2T-OUT-X312-LSmitll_OR2T-IN 0 z0=5 td=0.9ps
X295 X255-LSmitll_NDROT-OUT-X295-LSmitll_AND2T-IN X133-LSmitll_SPLITT-OUT-X295-LSmitll_AND2T-IN X486-LSmitll_SPLITT-OUT-X295-LSmitll_AND2T-IN X295-LSmitll_AND2T-OUT-X312-LSmitll_OR2T-INt LSmitll_AND2T

t1288 X296-LSmitll_AND2T-OUT-X312-LSmitll_OR2T-INt 0 X296-LSmitll_AND2T-OUT-X312-LSmitll_OR2T-IN 0 z0=5 td=9.2ps
X296 X131-LSmitll_SPLITT-OUT-X296-LSmitll_AND2T-IN X269-LSmitll_NDROT-OUT-X296-LSmitll_AND2T-IN X410-LSmitll_SPLITT-OUT-X296-LSmitll_AND2T-IN X296-LSmitll_AND2T-OUT-X312-LSmitll_OR2T-INt LSmitll_AND2T

t1289 X297-LSmitll_AND2T-OUT-X313-LSmitll_OR2T-INt 0 X297-LSmitll_AND2T-OUT-X313-LSmitll_OR2T-IN 0 z0=5 td=2.5ps
X297 X136-LSmitll_SPLITT-OUT-X297-LSmitll_AND2T-IN X229-LSmitll_NDROT-OUT-X297-LSmitll_AND2T-IN X568-LSmitll_SPLITT-OUT-X297-LSmitll_AND2T-IN X297-LSmitll_AND2T-OUT-X313-LSmitll_OR2T-INt LSmitll_AND2T

t1290 X298-LSmitll_AND2T-OUT-X313-LSmitll_OR2T-INt 0 X298-LSmitll_AND2T-OUT-X313-LSmitll_OR2T-IN 0 z0=5 td=19.2ps
X298 X123-LSmitll_SPLITT-OUT-X298-LSmitll_AND2T-IN X243-LSmitll_NDROT-OUT-X298-LSmitll_AND2T-IN X489-LSmitll_SPLITT-OUT-X298-LSmitll_AND2T-IN X298-LSmitll_AND2T-OUT-X313-LSmitll_OR2T-INt LSmitll_AND2T

t1291 X299-LSmitll_AND2T-OUT-X314-LSmitll_OR2T-INt 0 X299-LSmitll_AND2T-OUT-X314-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X299 X133-LSmitll_SPLITT-OUT-X299-LSmitll_AND2T-IN X257-LSmitll_NDROT-OUT-X299-LSmitll_AND2T-IN X502-LSmitll_SPLITT-OUT-X299-LSmitll_AND2T-IN X299-LSmitll_AND2T-OUT-X314-LSmitll_OR2T-INt LSmitll_AND2T

t1292 X300-LSmitll_AND2T-OUT-X314-LSmitll_OR2T-INt 0 X300-LSmitll_AND2T-OUT-X314-LSmitll_OR2T-IN 0 z0=5 td=22.3ps
X300 X121-LSmitll_SPLITT-OUT-X300-LSmitll_AND2T-IN X271-LSmitll_NDROT-OUT-X300-LSmitll_AND2T-IN X381-LSmitll_SPLITT-OUT-X300-LSmitll_AND2T-IN X300-LSmitll_AND2T-OUT-X314-LSmitll_OR2T-INt LSmitll_AND2T

t1293 X301-LSmitll_OR2T-OUT-X315-LSmitll_OR2T-INt 0 X301-LSmitll_OR2T-OUT-X315-LSmitll_OR2T-IN 0 z0=5 td=6.4ps
X301 X273-LSmitll_AND2T-OUT-X301-LSmitll_OR2T-IN X274-LSmitll_AND2T-OUT-X301-LSmitll_OR2T-IN X569-LSmitll_SPLITT-OUT-X301-LSmitll_OR2T-IN X301-LSmitll_OR2T-OUT-X315-LSmitll_OR2T-INt LSmitll_OR2T

t1294 X302-LSmitll_OR2T-OUT-X315-LSmitll_OR2T-INt 0 X302-LSmitll_OR2T-OUT-X315-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X302 X275-LSmitll_AND2T-OUT-X302-LSmitll_OR2T-IN X276-LSmitll_AND2T-OUT-X302-LSmitll_OR2T-IN X348-LSmitll_SPLITT-OUT-X302-LSmitll_OR2T-IN X302-LSmitll_OR2T-OUT-X315-LSmitll_OR2T-INt LSmitll_OR2T

t1295 X303-LSmitll_OR2T-OUT-X316-LSmitll_OR2T-INt 0 X303-LSmitll_OR2T-OUT-X316-LSmitll_OR2T-IN 0 z0=5 td=18.8ps
X303 X277-LSmitll_AND2T-OUT-X303-LSmitll_OR2T-IN X278-LSmitll_AND2T-OUT-X303-LSmitll_OR2T-IN X570-LSmitll_SPLITT-OUT-X303-LSmitll_OR2T-IN X303-LSmitll_OR2T-OUT-X316-LSmitll_OR2T-INt LSmitll_OR2T

t1296 X304-LSmitll_OR2T-OUT-X316-LSmitll_OR2T-INt 0 X304-LSmitll_OR2T-OUT-X316-LSmitll_OR2T-IN 0 z0=5 td=2.6ps
X304 X279-LSmitll_AND2T-OUT-X304-LSmitll_OR2T-IN X280-LSmitll_AND2T-OUT-X304-LSmitll_OR2T-IN X330-LSmitll_SPLITT-OUT-X304-LSmitll_OR2T-IN X304-LSmitll_OR2T-OUT-X316-LSmitll_OR2T-INt LSmitll_OR2T

t1297 X305-LSmitll_OR2T-OUT-X317-LSmitll_OR2T-INt 0 X305-LSmitll_OR2T-OUT-X317-LSmitll_OR2T-IN 0 z0=5 td=6.5ps
X305 X281-LSmitll_AND2T-OUT-X305-LSmitll_OR2T-IN X282-LSmitll_AND2T-OUT-X305-LSmitll_OR2T-IN X436-LSmitll_SPLITT-OUT-X305-LSmitll_OR2T-IN X305-LSmitll_OR2T-OUT-X317-LSmitll_OR2T-INt LSmitll_OR2T

t1298 X306-LSmitll_OR2T-OUT-X317-LSmitll_OR2T-INt 0 X306-LSmitll_OR2T-OUT-X317-LSmitll_OR2T-IN 0 z0=5 td=2.7ps
X306 X283-LSmitll_AND2T-OUT-X306-LSmitll_OR2T-IN X284-LSmitll_AND2T-OUT-X306-LSmitll_OR2T-IN X571-LSmitll_SPLITT-OUT-X306-LSmitll_OR2T-IN X306-LSmitll_OR2T-OUT-X317-LSmitll_OR2T-INt LSmitll_OR2T

t1299 X307-LSmitll_OR2T-OUT-X318-LSmitll_OR2T-INt 0 X307-LSmitll_OR2T-OUT-X318-LSmitll_OR2T-IN 0 z0=5 td=1.1ps
X307 X285-LSmitll_AND2T-OUT-X307-LSmitll_OR2T-IN X286-LSmitll_AND2T-OUT-X307-LSmitll_OR2T-IN X475-LSmitll_SPLITT-OUT-X307-LSmitll_OR2T-IN X307-LSmitll_OR2T-OUT-X318-LSmitll_OR2T-INt LSmitll_OR2T

t1300 X308-LSmitll_OR2T-OUT-X318-LSmitll_OR2T-INt 0 X308-LSmitll_OR2T-OUT-X318-LSmitll_OR2T-IN 0 z0=5 td=2.3ps
X308 X287-LSmitll_AND2T-OUT-X308-LSmitll_OR2T-IN X288-LSmitll_AND2T-OUT-X308-LSmitll_OR2T-IN X439-LSmitll_SPLITT-OUT-X308-LSmitll_OR2T-IN X308-LSmitll_OR2T-OUT-X318-LSmitll_OR2T-INt LSmitll_OR2T

t1301 X309-LSmitll_OR2T-OUT-X319-LSmitll_OR2T-INt 0 X309-LSmitll_OR2T-OUT-X319-LSmitll_OR2T-IN 0 z0=5 td=0.9ps
X309 X289-LSmitll_AND2T-OUT-X309-LSmitll_OR2T-IN X290-LSmitll_AND2T-OUT-X309-LSmitll_OR2T-IN X406-LSmitll_SPLITT-OUT-X309-LSmitll_OR2T-IN X309-LSmitll_OR2T-OUT-X319-LSmitll_OR2T-INt LSmitll_OR2T

t1302 X310-LSmitll_OR2T-OUT-X319-LSmitll_OR2T-INt 0 X310-LSmitll_OR2T-OUT-X319-LSmitll_OR2T-IN 0 z0=5 td=4.0ps
X310 X291-LSmitll_AND2T-OUT-X310-LSmitll_OR2T-IN X292-LSmitll_AND2T-OUT-X310-LSmitll_OR2T-IN X572-LSmitll_SPLITT-OUT-X310-LSmitll_OR2T-IN X310-LSmitll_OR2T-OUT-X319-LSmitll_OR2T-INt LSmitll_OR2T

t1303 X311-LSmitll_OR2T-OUT-X320-LSmitll_OR2T-INt 0 X311-LSmitll_OR2T-OUT-X320-LSmitll_OR2T-IN 0 z0=5 td=9.2ps
X311 X293-LSmitll_AND2T-OUT-X311-LSmitll_OR2T-IN X294-LSmitll_AND2T-OUT-X311-LSmitll_OR2T-IN X486-LSmitll_SPLITT-OUT-X311-LSmitll_OR2T-IN X311-LSmitll_OR2T-OUT-X320-LSmitll_OR2T-INt LSmitll_OR2T

t1304 X312-LSmitll_OR2T-OUT-X320-LSmitll_OR2T-INt 0 X312-LSmitll_OR2T-OUT-X320-LSmitll_OR2T-IN 0 z0=5 td=4.5ps
X312 X295-LSmitll_AND2T-OUT-X312-LSmitll_OR2T-IN X296-LSmitll_AND2T-OUT-X312-LSmitll_OR2T-IN X573-LSmitll_SPLITT-OUT-X312-LSmitll_OR2T-IN X312-LSmitll_OR2T-OUT-X320-LSmitll_OR2T-INt LSmitll_OR2T

t1305 X313-LSmitll_OR2T-OUT-X321-LSmitll_OR2T-INt 0 X313-LSmitll_OR2T-OUT-X321-LSmitll_OR2T-IN 0 z0=5 td=23.7ps
X313 X297-LSmitll_AND2T-OUT-X313-LSmitll_OR2T-IN X298-LSmitll_AND2T-OUT-X313-LSmitll_OR2T-IN X415-LSmitll_SPLITT-OUT-X313-LSmitll_OR2T-IN X313-LSmitll_OR2T-OUT-X321-LSmitll_OR2T-INt LSmitll_OR2T

t1306 X314-LSmitll_OR2T-OUT-X321-LSmitll_OR2T-INt 0 X314-LSmitll_OR2T-OUT-X321-LSmitll_OR2T-IN 0 z0=5 td=2.9ps
X314 X299-LSmitll_AND2T-OUT-X314-LSmitll_OR2T-IN X300-LSmitll_AND2T-OUT-X314-LSmitll_OR2T-IN X482-LSmitll_SPLITT-OUT-X314-LSmitll_OR2T-IN X314-LSmitll_OR2T-OUT-X321-LSmitll_OR2T-INt LSmitll_OR2T


X315 X301-LSmitll_OR2T-OUT-X315-LSmitll_OR2T-IN X302-LSmitll_OR2T-OUT-X315-LSmitll_OR2T-IN X574-LSmitll_SPLITT-OUT-X315-LSmitll_OR2T-IN bit_out0t LSmitll_OR2T


X316 X303-LSmitll_OR2T-OUT-X316-LSmitll_OR2T-IN X304-LSmitll_OR2T-OUT-X316-LSmitll_OR2T-IN X335-LSmitll_SPLITT-OUT-X316-LSmitll_OR2T-IN bit_out1t LSmitll_OR2T


X317 X305-LSmitll_OR2T-OUT-X317-LSmitll_OR2T-IN X306-LSmitll_OR2T-OUT-X317-LSmitll_OR2T-IN X362-LSmitll_SPLITT-OUT-X317-LSmitll_OR2T-IN bit_out2t LSmitll_OR2T


X318 X307-LSmitll_OR2T-OUT-X318-LSmitll_OR2T-IN X308-LSmitll_OR2T-OUT-X318-LSmitll_OR2T-IN X475-LSmitll_SPLITT-OUT-X318-LSmitll_OR2T-IN bit_out3t LSmitll_OR2T


X319 X309-LSmitll_OR2T-OUT-X319-LSmitll_OR2T-IN X310-LSmitll_OR2T-OUT-X319-LSmitll_OR2T-IN X410-LSmitll_SPLITT-OUT-X319-LSmitll_OR2T-IN bit_out4t LSmitll_OR2T


X320 X311-LSmitll_OR2T-OUT-X320-LSmitll_OR2T-IN X312-LSmitll_OR2T-OUT-X320-LSmitll_OR2T-IN X575-LSmitll_SPLITT-OUT-X320-LSmitll_OR2T-IN bit_out5t LSmitll_OR2T


X321 X313-LSmitll_OR2T-OUT-X321-LSmitll_OR2T-IN X314-LSmitll_OR2T-OUT-X321-LSmitll_OR2T-IN X492-LSmitll_SPLITT-OUT-X321-LSmitll_OR2T-IN bit_out6t LSmitll_OR2T

t1314 X322-LSmitll_SPLITT-OUT-X261-LSmitll_NDROT-INt 0 X322-LSmitll_SPLITT-OUT-X261-LSmitll_NDROT-IN 0 z0=5 td=2.8ps
t1315 X322-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-INt 0 X322-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X322 X324-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-IN X322-LSmitll_SPLITT-OUT-X261-LSmitll_NDROT-INt X322-LSmitll_SPLITT-OUT-X262-LSmitll_AND2T-INt LSmitll_SPLITT

t1316 X323-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-INt 0 X323-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-IN 0 z0=5 td=1.7ps
t1317 X323-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-INt 0 X323-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X323 X324-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-IN X323-LSmitll_SPLITT-OUT-X26-LSmitll_DFFT-INt X323-LSmitll_SPLITT-OUT-X28-LSmitll_DFFT-INt LSmitll_SPLITT

t1318 X324-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-INt 0 X324-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1319 X324-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-INt 0 X324-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X324 X327-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-IN X324-LSmitll_SPLITT-OUT-X322-LSmitll_SPLITT-INt X324-LSmitll_SPLITT-OUT-X323-LSmitll_SPLITT-INt LSmitll_SPLITT

t1320 X325-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-INt 0 X325-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1321 X325-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-INt 0 X325-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
X325 X326-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-IN X325-LSmitll_SPLITT-OUT-X63-LSmitll_DFFT-INt X325-LSmitll_SPLITT-OUT-X64-LSmitll_DFFT-INt LSmitll_SPLITT

t1322 X326-LSmitll_SPLITT-OUT-X566-LSmitll_SPLITT-INt 0 X326-LSmitll_SPLITT-OUT-X566-LSmitll_SPLITT-IN 0 z0=5 td=3.2ps
t1323 X326-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-INt 0 X326-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X326 X327-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-IN X326-LSmitll_SPLITT-OUT-X566-LSmitll_SPLITT-INt X326-LSmitll_SPLITT-OUT-X325-LSmitll_SPLITT-INt LSmitll_SPLITT

t1324 X327-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-INt 0 X327-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1325 X327-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-INt 0 X327-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X327 X333-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-IN X327-LSmitll_SPLITT-OUT-X324-LSmitll_SPLITT-INt X327-LSmitll_SPLITT-OUT-X326-LSmitll_SPLITT-INt LSmitll_SPLITT

t1326 X328-LSmitll_SPLITT-OUT-X27-LSmitll_DFFT-INt 0 X328-LSmitll_SPLITT-OUT-X27-LSmitll_DFFT-IN 0 z0=5 td=1.7ps
t1327 X328-LSmitll_SPLITT-OUT-X276-LSmitll_AND2T-INt 0 X328-LSmitll_SPLITT-OUT-X276-LSmitll_AND2T-IN 0 z0=5 td=0.5ps
X328 X329-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-IN X328-LSmitll_SPLITT-OUT-X27-LSmitll_DFFT-INt X328-LSmitll_SPLITT-OUT-X276-LSmitll_AND2T-INt LSmitll_SPLITT

t1328 X329-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-INt 0 X329-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-IN 0 z0=5 td=3.4ps
t1329 X329-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-INt 0 X329-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
X329 X332-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-IN X329-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-INt X329-LSmitll_SPLITT-OUT-X328-LSmitll_SPLITT-INt LSmitll_SPLITT

t1330 X330-LSmitll_SPLITT-OUT-X247-LSmitll_NDROT-INt 0 X330-LSmitll_SPLITT-OUT-X247-LSmitll_NDROT-IN 0 z0=5 td=2.6ps
t1331 X330-LSmitll_SPLITT-OUT-X304-LSmitll_OR2T-INt 0 X330-LSmitll_SPLITT-OUT-X304-LSmitll_OR2T-IN 0 z0=5 td=1.4ps
X330 X331-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-IN X330-LSmitll_SPLITT-OUT-X247-LSmitll_NDROT-INt X330-LSmitll_SPLITT-OUT-X304-LSmitll_OR2T-INt LSmitll_SPLITT

t1332 X331-LSmitll_SPLITT-OUT-X567-LSmitll_SPLITT-INt 0 X331-LSmitll_SPLITT-OUT-X567-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1333 X331-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-INt 0 X331-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X331 X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-IN X331-LSmitll_SPLITT-OUT-X567-LSmitll_SPLITT-INt X331-LSmitll_SPLITT-OUT-X330-LSmitll_SPLITT-INt LSmitll_SPLITT

t1334 X332-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-INt 0 X332-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1335 X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-INt 0 X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X332 X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-IN X332-LSmitll_SPLITT-OUT-X329-LSmitll_SPLITT-INt X332-LSmitll_SPLITT-OUT-X331-LSmitll_SPLITT-INt LSmitll_SPLITT

t1336 X333-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-INt 0 X333-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1337 X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-INt 0 X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-IN 0 z0=5 td=2.8ps
X333 X346-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-IN X333-LSmitll_SPLITT-OUT-X327-LSmitll_SPLITT-INt X333-LSmitll_SPLITT-OUT-X332-LSmitll_SPLITT-INt LSmitll_SPLITT

t1338 X334-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-INt 0 X334-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t1339 X334-LSmitll_SPLITT-OUT-X100-LSmitll_DFFT-INt 0 X334-LSmitll_SPLITT-OUT-X100-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
X334 X336-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-IN X334-LSmitll_SPLITT-OUT-X62-LSmitll_DFFT-INt X334-LSmitll_SPLITT-OUT-X100-LSmitll_DFFT-INt LSmitll_SPLITT

t1340 X335-LSmitll_SPLITT-OUT-X99-LSmitll_DFFT-INt 0 X335-LSmitll_SPLITT-OUT-X99-LSmitll_DFFT-IN 0 z0=5 td=5.6ps
t1341 X335-LSmitll_SPLITT-OUT-X316-LSmitll_OR2T-INt 0 X335-LSmitll_SPLITT-OUT-X316-LSmitll_OR2T-IN 0 z0=5 td=4.3ps
X335 X336-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-IN X335-LSmitll_SPLITT-OUT-X99-LSmitll_DFFT-INt X335-LSmitll_SPLITT-OUT-X316-LSmitll_OR2T-INt LSmitll_SPLITT

t1342 X336-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-INt 0 X336-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1343 X336-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-INt 0 X336-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X336 X339-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-IN X336-LSmitll_SPLITT-OUT-X334-LSmitll_SPLITT-INt X336-LSmitll_SPLITT-OUT-X335-LSmitll_SPLITT-INt LSmitll_SPLITT

t1344 X337-LSmitll_SPLITT-OUT-X98-LSmitll_DFFT-INt 0 X337-LSmitll_SPLITT-OUT-X98-LSmitll_DFFT-IN 0 z0=5 td=3.2ps
t1345 X337-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-INt 0 X337-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-IN 0 z0=5 td=1.8ps
X337 X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-IN X337-LSmitll_SPLITT-OUT-X98-LSmitll_DFFT-INt X337-LSmitll_SPLITT-OUT-X147-LSmitll_DFFT-INt LSmitll_SPLITT

t1346 X338-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-INt 0 X338-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1347 X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-INt 0 X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X338 X339-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-IN X338-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-INt X338-LSmitll_SPLITT-OUT-X337-LSmitll_SPLITT-INt LSmitll_SPLITT

t1348 X339-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-INt 0 X339-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-IN 0 z0=5 td=0.5ps
t1349 X339-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-INt 0 X339-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-IN 0 z0=5 td=3.7ps
X339 X345-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-IN X339-LSmitll_SPLITT-OUT-X336-LSmitll_SPLITT-INt X339-LSmitll_SPLITT-OUT-X338-LSmitll_SPLITT-INt LSmitll_SPLITT

t1350 X340-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-INt 0 X340-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-IN 0 z0=5 td=0.4ps
t1351 X340-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-INt 0 X340-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-IN 0 z0=5 td=3.2ps
X340 X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-IN X340-LSmitll_SPLITT-OUT-X264-LSmitll_AND2T-INt X340-LSmitll_SPLITT-OUT-X284-LSmitll_AND2T-INt LSmitll_SPLITT

t1352 X341-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-INt 0 X341-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1353 X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-INt 0 X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X341 X344-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-IN X341-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-INt X341-LSmitll_SPLITT-OUT-X340-LSmitll_SPLITT-INt LSmitll_SPLITT

t1354 X342-LSmitll_SPLITT-OUT-X265-LSmitll_NDROT-INt 0 X342-LSmitll_SPLITT-OUT-X265-LSmitll_NDROT-IN 0 z0=5 td=0.3ps
t1355 X342-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt 0 X342-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X342 X343-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-IN X342-LSmitll_SPLITT-OUT-X265-LSmitll_NDROT-INt X342-LSmitll_SPLITT-OUT-X266-LSmitll_AND2T-INt LSmitll_SPLITT

t1356 X343-LSmitll_SPLITT-OUT-X571-LSmitll_SPLITT-INt 0 X343-LSmitll_SPLITT-OUT-X571-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1357 X343-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-INt 0 X343-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
X343 X344-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-IN X343-LSmitll_SPLITT-OUT-X571-LSmitll_SPLITT-INt X343-LSmitll_SPLITT-OUT-X342-LSmitll_SPLITT-INt LSmitll_SPLITT

t1358 X344-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-INt 0 X344-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1359 X344-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-INt 0 X344-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X344 X345-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-IN X344-LSmitll_SPLITT-OUT-X341-LSmitll_SPLITT-INt X344-LSmitll_SPLITT-OUT-X343-LSmitll_SPLITT-INt LSmitll_SPLITT

t1360 X345-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-INt 0 X345-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1361 X345-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-INt 0 X345-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-IN 0 z0=5 td=3.7ps
X345 X346-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-IN X345-LSmitll_SPLITT-OUT-X339-LSmitll_SPLITT-INt X345-LSmitll_SPLITT-OUT-X344-LSmitll_SPLITT-INt LSmitll_SPLITT

t1362 X346-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-INt 0 X346-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-IN 0 z0=5 td=4.9ps
t1363 X346-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-INt 0 X346-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X346 X372-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-IN X346-LSmitll_SPLITT-OUT-X333-LSmitll_SPLITT-INt X346-LSmitll_SPLITT-OUT-X345-LSmitll_SPLITT-INt LSmitll_SPLITT

t1364 X347-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-INt 0 X347-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-IN 0 z0=5 td=1.5ps
t1365 X347-LSmitll_SPLITT-OUT-X259-LSmitll_NDROT-INt 0 X347-LSmitll_SPLITT-OUT-X259-LSmitll_NDROT-IN 0 z0=5 td=2.1ps
X347 X349-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-IN X347-LSmitll_SPLITT-OUT-X248-LSmitll_AND2T-INt X347-LSmitll_SPLITT-OUT-X259-LSmitll_NDROT-INt LSmitll_SPLITT

t1366 X348-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-INt 0 X348-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-IN 0 z0=5 td=2.0ps
t1367 X348-LSmitll_SPLITT-OUT-X302-LSmitll_OR2T-INt 0 X348-LSmitll_SPLITT-OUT-X302-LSmitll_OR2T-IN 0 z0=5 td=1.4ps
X348 X349-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-IN X348-LSmitll_SPLITT-OUT-X24-LSmitll_DFFT-INt X348-LSmitll_SPLITT-OUT-X302-LSmitll_OR2T-INt LSmitll_SPLITT

t1368 X349-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-INt 0 X349-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1369 X349-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-INt 0 X349-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X349 X352-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-IN X349-LSmitll_SPLITT-OUT-X347-LSmitll_SPLITT-INt X349-LSmitll_SPLITT-OUT-X348-LSmitll_SPLITT-INt LSmitll_SPLITT

t1370 X350-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-INt 0 X350-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t1371 X350-LSmitll_SPLITT-OUT-X279-LSmitll_AND2T-INt 0 X350-LSmitll_SPLITT-OUT-X279-LSmitll_AND2T-IN 0 z0=5 td=1.3ps
X350 X351-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-IN X350-LSmitll_SPLITT-OUT-X60-LSmitll_DFFT-INt X350-LSmitll_SPLITT-OUT-X279-LSmitll_AND2T-INt LSmitll_SPLITT

t1372 X351-LSmitll_SPLITT-OUT-X574-LSmitll_SPLITT-INt 0 X351-LSmitll_SPLITT-OUT-X574-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
t1373 X351-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-INt 0 X351-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X351 X352-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-IN X351-LSmitll_SPLITT-OUT-X574-LSmitll_SPLITT-INt X351-LSmitll_SPLITT-OUT-X350-LSmitll_SPLITT-INt LSmitll_SPLITT

t1374 X352-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-INt 0 X352-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1375 X352-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-INt 0 X352-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X352 X358-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-IN X352-LSmitll_SPLITT-OUT-X349-LSmitll_SPLITT-INt X352-LSmitll_SPLITT-OUT-X351-LSmitll_SPLITT-INt LSmitll_SPLITT

t1376 X353-LSmitll_SPLITT-OUT-X25-LSmitll_DFFT-INt 0 X353-LSmitll_SPLITT-OUT-X25-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
t1377 X353-LSmitll_SPLITT-OUT-X275-LSmitll_AND2T-INt 0 X353-LSmitll_SPLITT-OUT-X275-LSmitll_AND2T-IN 0 z0=5 td=0.8ps
X353 X354-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-IN X353-LSmitll_SPLITT-OUT-X25-LSmitll_DFFT-INt X353-LSmitll_SPLITT-OUT-X275-LSmitll_AND2T-INt LSmitll_SPLITT

t1378 X354-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-INt 0 X354-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1379 X354-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-INt 0 X354-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X354 X357-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-IN X354-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-INt X354-LSmitll_SPLITT-OUT-X353-LSmitll_SPLITT-INt LSmitll_SPLITT

t1380 X355-LSmitll_SPLITT-OUT-X233-LSmitll_NDROT-INt 0 X355-LSmitll_SPLITT-OUT-X233-LSmitll_NDROT-IN 0 z0=5 td=0.8ps
t1381 X355-LSmitll_SPLITT-OUT-X278-LSmitll_AND2T-INt 0 X355-LSmitll_SPLITT-OUT-X278-LSmitll_AND2T-IN 0 z0=5 td=0.5ps
X355 X356-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-IN X355-LSmitll_SPLITT-OUT-X233-LSmitll_NDROT-INt X355-LSmitll_SPLITT-OUT-X278-LSmitll_AND2T-INt LSmitll_SPLITT

t1382 X356-LSmitll_SPLITT-OUT-X569-LSmitll_SPLITT-INt 0 X356-LSmitll_SPLITT-OUT-X569-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
t1383 X356-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-INt 0 X356-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X356 X357-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-IN X356-LSmitll_SPLITT-OUT-X569-LSmitll_SPLITT-INt X356-LSmitll_SPLITT-OUT-X355-LSmitll_SPLITT-INt LSmitll_SPLITT

t1384 X357-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-INt 0 X357-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1385 X357-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-INt 0 X357-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X357 X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-IN X357-LSmitll_SPLITT-OUT-X354-LSmitll_SPLITT-INt X357-LSmitll_SPLITT-OUT-X356-LSmitll_SPLITT-INt LSmitll_SPLITT

t1386 X358-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-INt 0 X358-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1387 X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-INt 0 X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
X358 X371-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-IN X358-LSmitll_SPLITT-OUT-X352-LSmitll_SPLITT-INt X358-LSmitll_SPLITT-OUT-X357-LSmitll_SPLITT-INt LSmitll_SPLITT

t1388 X359-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-INt 0 X359-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t1389 X359-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt 0 X359-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-IN 0 z0=5 td=3.3ps
X359 X361-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-IN X359-LSmitll_SPLITT-OUT-X61-LSmitll_DFFT-INt X359-LSmitll_SPLITT-OUT-X101-LSmitll_AND2T-INt LSmitll_SPLITT

t1390 X360-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-INt 0 X360-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-IN 0 z0=5 td=0.5ps
t1391 X360-LSmitll_SPLITT-OUT-X249-LSmitll_NDROT-INt 0 X360-LSmitll_SPLITT-OUT-X249-LSmitll_NDROT-IN 0 z0=5 td=2.8ps
X360 X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-IN X360-LSmitll_SPLITT-OUT-X102-LSmitll_AND2T-INt X360-LSmitll_SPLITT-OUT-X249-LSmitll_NDROT-INt LSmitll_SPLITT

t1392 X361-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-INt 0 X361-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
t1393 X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-INt 0 X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X361 X364-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-IN X361-LSmitll_SPLITT-OUT-X359-LSmitll_SPLITT-INt X361-LSmitll_SPLITT-OUT-X360-LSmitll_SPLITT-INt LSmitll_SPLITT

t1394 X362-LSmitll_SPLITT-OUT-X288-LSmitll_AND2T-INt 0 X362-LSmitll_SPLITT-OUT-X288-LSmitll_AND2T-IN 0 z0=5 td=0.4ps
t1395 X362-LSmitll_SPLITT-OUT-X317-LSmitll_OR2T-INt 0 X362-LSmitll_SPLITT-OUT-X317-LSmitll_OR2T-IN 0 z0=5 td=1.7ps
X362 X363-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-IN X362-LSmitll_SPLITT-OUT-X288-LSmitll_AND2T-INt X362-LSmitll_SPLITT-OUT-X317-LSmitll_OR2T-INt LSmitll_SPLITT

t1396 X363-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-INt 0 X363-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1397 X363-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-INt 0 X363-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X363 X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-IN X363-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-INt X363-LSmitll_SPLITT-OUT-X362-LSmitll_SPLITT-INt LSmitll_SPLITT

t1398 X364-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-INt 0 X364-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1399 X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-INt 0 X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X364 X370-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-IN X364-LSmitll_SPLITT-OUT-X361-LSmitll_SPLITT-INt X364-LSmitll_SPLITT-OUT-X363-LSmitll_SPLITT-INt LSmitll_SPLITT

t1400 X365-LSmitll_SPLITT-OUT-X65-LSmitll_AND2T-INt 0 X365-LSmitll_SPLITT-OUT-X65-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1401 X365-LSmitll_SPLITT-OUT-X96-LSmitll_DFFT-INt 0 X365-LSmitll_SPLITT-OUT-X96-LSmitll_DFFT-IN 0 z0=5 td=0.3ps
X365 X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-IN X365-LSmitll_SPLITT-OUT-X65-LSmitll_AND2T-INt X365-LSmitll_SPLITT-OUT-X96-LSmitll_DFFT-INt LSmitll_SPLITT

t1402 X366-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-INt 0 X366-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1403 X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-INt 0 X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X366 X369-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-IN X366-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-INt X366-LSmitll_SPLITT-OUT-X365-LSmitll_SPLITT-INt LSmitll_SPLITT

t1404 X367-LSmitll_SPLITT-OUT-X95-LSmitll_DFFT-INt 0 X367-LSmitll_SPLITT-OUT-X95-LSmitll_DFFT-IN 0 z0=5 td=11.3ps
t1405 X367-LSmitll_SPLITT-OUT-X251-LSmitll_NDROT-INt 0 X367-LSmitll_SPLITT-OUT-X251-LSmitll_NDROT-IN 0 z0=5 td=1.0ps
X367 X368-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-IN X367-LSmitll_SPLITT-OUT-X95-LSmitll_DFFT-INt X367-LSmitll_SPLITT-OUT-X251-LSmitll_NDROT-INt LSmitll_SPLITT

t1406 X368-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-INt 0 X368-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1407 X368-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-INt 0 X368-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X368 X369-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-IN X368-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-INt X368-LSmitll_SPLITT-OUT-X367-LSmitll_SPLITT-INt LSmitll_SPLITT

t1408 X369-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-INt 0 X369-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
t1409 X369-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-INt 0 X369-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X369 X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-IN X369-LSmitll_SPLITT-OUT-X366-LSmitll_SPLITT-INt X369-LSmitll_SPLITT-OUT-X368-LSmitll_SPLITT-INt LSmitll_SPLITT

t1410 X370-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-INt 0 X370-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t1411 X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-INt 0 X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-IN 0 z0=5 td=3.5ps
X370 X371-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-IN X370-LSmitll_SPLITT-OUT-X364-LSmitll_SPLITT-INt X370-LSmitll_SPLITT-OUT-X369-LSmitll_SPLITT-INt LSmitll_SPLITT

t1412 X371-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-INt 0 X371-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1413 X371-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-INt 0 X371-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-IN 0 z0=5 td=4.7ps
X371 X372-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-IN X371-LSmitll_SPLITT-OUT-X358-LSmitll_SPLITT-INt X371-LSmitll_SPLITT-OUT-X370-LSmitll_SPLITT-INt LSmitll_SPLITT

t1414 X372-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-INt 0 X372-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-IN 0 z0=5 td=4.7ps
t1415 X372-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-INt 0 X372-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-IN 0 z0=5 td=4.3ps
X372 X423-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-IN X372-LSmitll_SPLITT-OUT-X346-LSmitll_SPLITT-INt X372-LSmitll_SPLITT-OUT-X371-LSmitll_SPLITT-INt LSmitll_SPLITT

t1416 X373-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-INt 0 X373-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
t1417 X373-LSmitll_SPLITT-OUT-X148-LSmitll_DFFT-INt 0 X373-LSmitll_SPLITT-OUT-X148-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
X373 X375-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-IN X373-LSmitll_SPLITT-OUT-X146-LSmitll_DFFT-INt X373-LSmitll_SPLITT-OUT-X148-LSmitll_DFFT-INt LSmitll_SPLITT

t1418 X374-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-INt 0 X374-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-IN 0 z0=5 td=3.8ps
t1419 X374-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-INt 0 X374-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
X374 X375-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-IN X374-LSmitll_SPLITT-OUT-X30-LSmitll_DFFT-INt X374-LSmitll_SPLITT-OUT-X167-LSmitll_DFFT-INt LSmitll_SPLITT

t1420 X375-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-INt 0 X375-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1421 X375-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-INt 0 X375-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X375 X378-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-IN X375-LSmitll_SPLITT-OUT-X373-LSmitll_SPLITT-INt X375-LSmitll_SPLITT-OUT-X374-LSmitll_SPLITT-INt LSmitll_SPLITT

t1422 X376-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-INt 0 X376-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-IN 0 z0=5 td=1.5ps
t1423 X376-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-INt 0 X376-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
X376 X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-IN X376-LSmitll_SPLITT-OUT-X186-LSmitll_DFFT-INt X376-LSmitll_SPLITT-OUT-X187-LSmitll_DFFT-INt LSmitll_SPLITT

t1424 X377-LSmitll_SPLITT-OUT-X564-LSmitll_SPLITT-INt 0 X377-LSmitll_SPLITT-OUT-X564-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1425 X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-INt 0 X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X377 X378-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-IN X377-LSmitll_SPLITT-OUT-X564-LSmitll_SPLITT-INt X377-LSmitll_SPLITT-OUT-X376-LSmitll_SPLITT-INt LSmitll_SPLITT

t1426 X378-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-INt 0 X378-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1427 X378-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-INt 0 X378-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X378 X384-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-IN X378-LSmitll_SPLITT-OUT-X375-LSmitll_SPLITT-INt X378-LSmitll_SPLITT-OUT-X377-LSmitll_SPLITT-INt LSmitll_SPLITT

t1428 X379-LSmitll_SPLITT-OUT-X67-LSmitll_AND2T-INt 0 X379-LSmitll_SPLITT-OUT-X67-LSmitll_AND2T-IN 0 z0=5 td=3.0ps
t1429 X379-LSmitll_SPLITT-OUT-X168-LSmitll_DFFT-INt 0 X379-LSmitll_SPLITT-OUT-X168-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
X379 X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-IN X379-LSmitll_SPLITT-OUT-X67-LSmitll_AND2T-INt X379-LSmitll_SPLITT-OUT-X168-LSmitll_DFFT-INt LSmitll_SPLITT

t1430 X380-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-INt 0 X380-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1431 X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-INt 0 X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X380 X383-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-IN X380-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-INt X380-LSmitll_SPLITT-OUT-X379-LSmitll_SPLITT-INt LSmitll_SPLITT

t1432 X381-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-INt 0 X381-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-IN 0 z0=5 td=0.8ps
t1433 X381-LSmitll_SPLITT-OUT-X300-LSmitll_AND2T-INt 0 X381-LSmitll_SPLITT-OUT-X300-LSmitll_AND2T-IN 0 z0=5 td=3.6ps
X381 X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-IN X381-LSmitll_SPLITT-OUT-X270-LSmitll_AND2T-INt X381-LSmitll_SPLITT-OUT-X300-LSmitll_AND2T-INt LSmitll_SPLITT

t1434 X382-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-INt 0 X382-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
t1435 X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-INt 0 X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X382 X383-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-IN X382-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-INt X382-LSmitll_SPLITT-OUT-X381-LSmitll_SPLITT-INt LSmitll_SPLITT

t1436 X383-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-INt 0 X383-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1437 X383-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-INt 0 X383-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X383 X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-IN X383-LSmitll_SPLITT-OUT-X380-LSmitll_SPLITT-INt X383-LSmitll_SPLITT-OUT-X382-LSmitll_SPLITT-INt LSmitll_SPLITT

t1438 X384-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-INt 0 X384-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1439 X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-INt 0 X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X384 X397-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-IN X384-LSmitll_SPLITT-OUT-X378-LSmitll_SPLITT-INt X384-LSmitll_SPLITT-OUT-X383-LSmitll_SPLITT-INt LSmitll_SPLITT

t1440 X385-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-INt 0 X385-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-IN 0 z0=5 td=5.0ps
t1441 X385-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-INt 0 X385-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
X385 X387-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-IN X385-LSmitll_SPLITT-OUT-X161-LSmitll_DFFT-INt X385-LSmitll_SPLITT-OUT-X188-LSmitll_DFFT-INt LSmitll_SPLITT

t1442 X386-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt 0 X386-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
t1443 X386-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-INt 0 X386-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-IN 0 z0=5 td=2.2ps
X386 X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-IN X386-LSmitll_SPLITT-OUT-X240-LSmitll_AND2T-INt X386-LSmitll_SPLITT-OUT-X272-LSmitll_AND2T-INt LSmitll_SPLITT

t1444 X387-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-INt 0 X387-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1445 X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-INt 0 X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
X387 X390-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-IN X387-LSmitll_SPLITT-OUT-X385-LSmitll_SPLITT-INt X387-LSmitll_SPLITT-OUT-X386-LSmitll_SPLITT-INt LSmitll_SPLITT

t1446 X388-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-INt 0 X388-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-IN 0 z0=5 td=4.0ps
t1447 X388-LSmitll_SPLITT-OUT-X162-LSmitll_DFFT-INt 0 X388-LSmitll_SPLITT-OUT-X162-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X388 X389-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-IN X388-LSmitll_SPLITT-OUT-X31-LSmitll_DFFT-INt X388-LSmitll_SPLITT-OUT-X162-LSmitll_DFFT-INt LSmitll_SPLITT

t1448 X389-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-INt 0 X389-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1449 X389-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-INt 0 X389-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X389 X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-IN X389-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-INt X389-LSmitll_SPLITT-OUT-X388-LSmitll_SPLITT-INt LSmitll_SPLITT

t1450 X390-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-INt 0 X390-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1451 X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-INt 0 X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
X390 X396-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-IN X390-LSmitll_SPLITT-OUT-X387-LSmitll_SPLITT-INt X390-LSmitll_SPLITT-OUT-X389-LSmitll_SPLITT-INt LSmitll_SPLITT

t1452 X391-LSmitll_SPLITT-OUT-X239-LSmitll_NDROT-INt 0 X391-LSmitll_SPLITT-OUT-X239-LSmitll_NDROT-IN 0 z0=5 td=2.7ps
t1453 X391-LSmitll_SPLITT-OUT-X290-LSmitll_AND2T-INt 0 X391-LSmitll_SPLITT-OUT-X290-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
X391 X392-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-IN X391-LSmitll_SPLITT-OUT-X239-LSmitll_NDROT-INt X391-LSmitll_SPLITT-OUT-X290-LSmitll_AND2T-INt LSmitll_SPLITT

t1454 X392-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-INt 0 X392-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1455 X392-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-INt 0 X392-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X392 X395-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-IN X392-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-INt X392-LSmitll_SPLITT-OUT-X391-LSmitll_SPLITT-INt LSmitll_SPLITT

t1456 X393-LSmitll_SPLITT-OUT-X39-LSmitll_NOTT-INt 0 X393-LSmitll_SPLITT-OUT-X39-LSmitll_NOTT-IN 0 z0=5 td=1.2ps
t1457 X393-LSmitll_SPLITT-OUT-X70-LSmitll_AND2T-INt 0 X393-LSmitll_SPLITT-OUT-X70-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
X393 X394-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-IN X393-LSmitll_SPLITT-OUT-X39-LSmitll_NOTT-INt X393-LSmitll_SPLITT-OUT-X70-LSmitll_AND2T-INt LSmitll_SPLITT

t1458 X394-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-INt 0 X394-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1459 X394-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-INt 0 X394-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X394 X395-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-IN X394-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-INt X394-LSmitll_SPLITT-OUT-X393-LSmitll_SPLITT-INt LSmitll_SPLITT

t1460 X395-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-INt 0 X395-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1461 X395-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-INt 0 X395-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X395 X396-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-IN X395-LSmitll_SPLITT-OUT-X392-LSmitll_SPLITT-INt X395-LSmitll_SPLITT-OUT-X394-LSmitll_SPLITT-INt LSmitll_SPLITT

t1462 X396-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-INt 0 X396-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1463 X396-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-INt 0 X396-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-IN 0 z0=5 td=3.4ps
X396 X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-IN X396-LSmitll_SPLITT-OUT-X390-LSmitll_SPLITT-INt X396-LSmitll_SPLITT-OUT-X395-LSmitll_SPLITT-INt LSmitll_SPLITT

t1464 X397-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-INt 0 X397-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-IN 0 z0=5 td=3.4ps
t1465 X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-INt 0 X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
X397 X422-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-IN X397-LSmitll_SPLITT-OUT-X384-LSmitll_SPLITT-INt X397-LSmitll_SPLITT-OUT-X396-LSmitll_SPLITT-INt LSmitll_SPLITT

t1466 X398-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-INt 0 X398-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-IN 0 z0=5 td=3.6ps
t1467 X398-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-INt 0 X398-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-IN 0 z0=5 td=0.3ps
X398 X400-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-IN X398-LSmitll_SPLITT-OUT-X144-LSmitll_DFFT-INt X398-LSmitll_SPLITT-OUT-X268-LSmitll_AND2T-INt LSmitll_SPLITT

t1468 X399-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-INt 0 X399-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-IN 0 z0=5 td=3.8ps
t1469 X399-LSmitll_SPLITT-OUT-X267-LSmitll_NDROT-INt 0 X399-LSmitll_SPLITT-OUT-X267-LSmitll_NDROT-IN 0 z0=5 td=0.5ps
X399 X400-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-IN X399-LSmitll_SPLITT-OUT-X145-LSmitll_DFFT-INt X399-LSmitll_SPLITT-OUT-X267-LSmitll_NDROT-INt LSmitll_SPLITT

t1470 X400-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-INt 0 X400-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1471 X400-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-INt 0 X400-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X400 X403-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-IN X400-LSmitll_SPLITT-OUT-X398-LSmitll_SPLITT-INt X400-LSmitll_SPLITT-OUT-X399-LSmitll_SPLITT-INt LSmitll_SPLITT

t1472 X401-LSmitll_SPLITT-OUT-X269-LSmitll_NDROT-INt 0 X401-LSmitll_SPLITT-OUT-X269-LSmitll_NDROT-IN 0 z0=5 td=1.7ps
t1473 X401-LSmitll_SPLITT-OUT-X292-LSmitll_AND2T-INt 0 X401-LSmitll_SPLITT-OUT-X292-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
X401 X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-IN X401-LSmitll_SPLITT-OUT-X269-LSmitll_NDROT-INt X401-LSmitll_SPLITT-OUT-X292-LSmitll_AND2T-INt LSmitll_SPLITT

t1474 X402-LSmitll_SPLITT-OUT-X572-LSmitll_SPLITT-INt 0 X402-LSmitll_SPLITT-OUT-X572-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1475 X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-INt 0 X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X402 X403-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-IN X402-LSmitll_SPLITT-OUT-X572-LSmitll_SPLITT-INt X402-LSmitll_SPLITT-OUT-X401-LSmitll_SPLITT-INt LSmitll_SPLITT

t1476 X403-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-INt 0 X403-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-IN 0 z0=5 td=0.5ps
t1477 X403-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-INt 0 X403-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X403 X409-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-IN X403-LSmitll_SPLITT-OUT-X400-LSmitll_SPLITT-INt X403-LSmitll_SPLITT-OUT-X402-LSmitll_SPLITT-INt LSmitll_SPLITT

t1478 X404-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-INt 0 X404-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
t1479 X404-LSmitll_SPLITT-OUT-X287-LSmitll_AND2T-INt 0 X404-LSmitll_SPLITT-OUT-X287-LSmitll_AND2T-IN 0 z0=5 td=0.7ps
X404 X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-IN X404-LSmitll_SPLITT-OUT-X143-LSmitll_DFFT-INt X404-LSmitll_SPLITT-OUT-X287-LSmitll_AND2T-INt LSmitll_SPLITT

t1480 X405-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-INt 0 X405-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1481 X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-INt 0 X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
X405 X408-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-IN X405-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-INt X405-LSmitll_SPLITT-OUT-X404-LSmitll_SPLITT-INt LSmitll_SPLITT

t1482 X406-LSmitll_SPLITT-OUT-X291-LSmitll_AND2T-INt 0 X406-LSmitll_SPLITT-OUT-X291-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
t1483 X406-LSmitll_SPLITT-OUT-X309-LSmitll_OR2T-INt 0 X406-LSmitll_SPLITT-OUT-X309-LSmitll_OR2T-IN 0 z0=5 td=3.4ps
X406 X407-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-IN X406-LSmitll_SPLITT-OUT-X291-LSmitll_AND2T-INt X406-LSmitll_SPLITT-OUT-X309-LSmitll_OR2T-INt LSmitll_SPLITT

t1484 X407-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-INt 0 X407-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-IN 0 z0=5 td=2.8ps
t1485 X407-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-INt 0 X407-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X407 X408-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-IN X407-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-INt X407-LSmitll_SPLITT-OUT-X406-LSmitll_SPLITT-INt LSmitll_SPLITT

t1486 X408-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-INt 0 X408-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1487 X408-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-INt 0 X408-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X408 X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-IN X408-LSmitll_SPLITT-OUT-X405-LSmitll_SPLITT-INt X408-LSmitll_SPLITT-OUT-X407-LSmitll_SPLITT-INt LSmitll_SPLITT

t1488 X409-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-INt 0 X409-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1489 X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-INt 0 X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X409 X421-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-IN X409-LSmitll_SPLITT-OUT-X403-LSmitll_SPLITT-INt X409-LSmitll_SPLITT-OUT-X408-LSmitll_SPLITT-INt LSmitll_SPLITT

t1490 X410-LSmitll_SPLITT-OUT-X296-LSmitll_AND2T-INt 0 X410-LSmitll_SPLITT-OUT-X296-LSmitll_AND2T-IN 0 z0=5 td=1.5ps
t1491 X410-LSmitll_SPLITT-OUT-X319-LSmitll_OR2T-INt 0 X410-LSmitll_SPLITT-OUT-X319-LSmitll_OR2T-IN 0 z0=5 td=1.3ps
X410 X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-IN X410-LSmitll_SPLITT-OUT-X296-LSmitll_AND2T-INt X410-LSmitll_SPLITT-OUT-X319-LSmitll_OR2T-INt LSmitll_SPLITT

t1492 X411-LSmitll_SPLITT-OUT-X568-LSmitll_SPLITT-INt 0 X411-LSmitll_SPLITT-OUT-X568-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
t1493 X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-INt 0 X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-IN 0 z0=5 td=0.5ps
X411 X414-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-IN X411-LSmitll_SPLITT-OUT-X568-LSmitll_SPLITT-INt X411-LSmitll_SPLITT-OUT-X410-LSmitll_SPLITT-INt LSmitll_SPLITT

t1494 X412-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-INt 0 X412-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-IN 0 z0=5 td=3.1ps
t1495 X412-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-INt 0 X412-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
X412 X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-IN X412-LSmitll_SPLITT-OUT-X34-LSmitll_OR2T-INt X412-LSmitll_SPLITT-OUT-X108-LSmitll_AND2T-INt LSmitll_SPLITT

t1496 X413-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-INt 0 X413-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1497 X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-INt 0 X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X413 X414-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-IN X413-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-INt X413-LSmitll_SPLITT-OUT-X412-LSmitll_SPLITT-INt LSmitll_SPLITT

t1498 X414-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-INt 0 X414-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1499 X414-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-INt 0 X414-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
X414 X420-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-IN X414-LSmitll_SPLITT-OUT-X411-LSmitll_SPLITT-INt X414-LSmitll_SPLITT-OUT-X413-LSmitll_SPLITT-INt LSmitll_SPLITT

t1500 X415-LSmitll_SPLITT-OUT-X293-LSmitll_AND2T-INt 0 X415-LSmitll_SPLITT-OUT-X293-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
t1501 X415-LSmitll_SPLITT-OUT-X313-LSmitll_OR2T-INt 0 X415-LSmitll_SPLITT-OUT-X313-LSmitll_OR2T-IN 0 z0=5 td=2.4ps
X415 X416-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-IN X415-LSmitll_SPLITT-OUT-X293-LSmitll_AND2T-INt X415-LSmitll_SPLITT-OUT-X313-LSmitll_OR2T-INt LSmitll_SPLITT

t1502 X416-LSmitll_SPLITT-OUT-X573-LSmitll_SPLITT-INt 0 X416-LSmitll_SPLITT-OUT-X573-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1503 X416-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-INt 0 X416-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
X416 X419-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-IN X416-LSmitll_SPLITT-OUT-X573-LSmitll_SPLITT-INt X416-LSmitll_SPLITT-OUT-X415-LSmitll_SPLITT-INt LSmitll_SPLITT

t1504 X417-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-INt 0 X417-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t1505 X417-LSmitll_SPLITT-OUT-X182-LSmitll_DFFT-INt 0 X417-LSmitll_SPLITT-OUT-X182-LSmitll_DFFT-IN 0 z0=5 td=1.2ps
X417 X418-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-IN X417-LSmitll_SPLITT-OUT-X181-LSmitll_DFFT-INt X417-LSmitll_SPLITT-OUT-X182-LSmitll_DFFT-INt LSmitll_SPLITT

t1506 X418-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-INt 0 X418-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1507 X418-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-INt 0 X418-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X418 X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-IN X418-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-INt X418-LSmitll_SPLITT-OUT-X417-LSmitll_SPLITT-INt LSmitll_SPLITT

t1508 X419-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-INt 0 X419-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1509 X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-INt 0 X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X419 X420-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-IN X419-LSmitll_SPLITT-OUT-X416-LSmitll_SPLITT-INt X419-LSmitll_SPLITT-OUT-X418-LSmitll_SPLITT-INt LSmitll_SPLITT

t1510 X420-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-INt 0 X420-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-IN 0 z0=5 td=2.8ps
t1511 X420-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-INt 0 X420-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X420 X421-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-IN X420-LSmitll_SPLITT-OUT-X414-LSmitll_SPLITT-INt X420-LSmitll_SPLITT-OUT-X419-LSmitll_SPLITT-INt LSmitll_SPLITT

t1512 X421-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-INt 0 X421-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-IN 0 z0=5 td=3.2ps
t1513 X421-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-INt 0 X421-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
X421 X422-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-IN X421-LSmitll_SPLITT-OUT-X409-LSmitll_SPLITT-INt X421-LSmitll_SPLITT-OUT-X420-LSmitll_SPLITT-INt LSmitll_SPLITT

t1514 X422-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-INt 0 X422-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-IN 0 z0=5 td=4.3ps
t1515 X422-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-INt 0 X422-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-IN 0 z0=5 td=5.5ps
X422 X423-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-IN X422-LSmitll_SPLITT-OUT-X397-LSmitll_SPLITT-INt X422-LSmitll_SPLITT-OUT-X421-LSmitll_SPLITT-INt LSmitll_SPLITT

t1516 X423-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-INt 0 X423-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-IN 0 z0=5 td=6.5ps
t1517 X423-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-INt 0 X423-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-IN 0 z0=5 td=3.5ps
X423 X576-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-IN X423-LSmitll_SPLITT-OUT-X372-LSmitll_SPLITT-INt X423-LSmitll_SPLITT-OUT-X422-LSmitll_SPLITT-INt LSmitll_SPLITT

t1518 X424-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-INt 0 X424-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-IN 0 z0=5 td=2.6ps
t1519 X424-LSmitll_SPLITT-OUT-X274-LSmitll_AND2T-INt 0 X424-LSmitll_SPLITT-OUT-X274-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
X424 X426-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-IN X424-LSmitll_SPLITT-OUT-X246-LSmitll_AND2T-INt X424-LSmitll_SPLITT-OUT-X274-LSmitll_AND2T-INt LSmitll_SPLITT

t1520 X425-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-INt 0 X425-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1521 X425-LSmitll_SPLITT-OUT-X231-LSmitll_NDROT-INt 0 X425-LSmitll_SPLITT-OUT-X231-LSmitll_NDROT-IN 0 z0=5 td=0.3ps
X425 X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-IN X425-LSmitll_SPLITT-OUT-X20-LSmitll_DFFT-INt X425-LSmitll_SPLITT-OUT-X231-LSmitll_NDROT-INt LSmitll_SPLITT

t1522 X426-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-INt 0 X426-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1523 X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-INt 0 X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X426 X429-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-IN X426-LSmitll_SPLITT-OUT-X424-LSmitll_SPLITT-INt X426-LSmitll_SPLITT-OUT-X425-LSmitll_SPLITT-INt LSmitll_SPLITT

t1524 X427-LSmitll_SPLITT-OUT-X37-LSmitll_NOTT-INt 0 X427-LSmitll_SPLITT-OUT-X37-LSmitll_NOTT-IN 0 z0=5 td=1.1ps
t1525 X427-LSmitll_SPLITT-OUT-X59-LSmitll_DFFT-INt 0 X427-LSmitll_SPLITT-OUT-X59-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
X427 X428-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-IN X427-LSmitll_SPLITT-OUT-X37-LSmitll_NOTT-INt X427-LSmitll_SPLITT-OUT-X59-LSmitll_DFFT-INt LSmitll_SPLITT

t1526 X428-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-INt 0 X428-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1527 X428-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-INt 0 X428-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-IN 0 z0=5 td=0.6ps
X428 X429-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-IN X428-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-INt X428-LSmitll_SPLITT-OUT-X427-LSmitll_SPLITT-INt LSmitll_SPLITT

t1528 X429-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-INt 0 X429-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1529 X429-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-INt 0 X429-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X429 X435-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-IN X429-LSmitll_SPLITT-OUT-X426-LSmitll_SPLITT-INt X429-LSmitll_SPLITT-OUT-X428-LSmitll_SPLITT-INt LSmitll_SPLITT

t1530 X430-LSmitll_SPLITT-OUT-X22-LSmitll_DFFT-INt 0 X430-LSmitll_SPLITT-OUT-X22-LSmitll_DFFT-IN 0 z0=5 td=2.1ps
t1531 X430-LSmitll_SPLITT-OUT-X23-LSmitll_DFFT-INt 0 X430-LSmitll_SPLITT-OUT-X23-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
X430 X431-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-IN X430-LSmitll_SPLITT-OUT-X22-LSmitll_DFFT-INt X430-LSmitll_SPLITT-OUT-X23-LSmitll_DFFT-INt LSmitll_SPLITT

t1532 X431-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-INt 0 X431-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1533 X431-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-INt 0 X431-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-IN 0 z0=5 td=0.6ps
X431 X434-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-IN X431-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-INt X431-LSmitll_SPLITT-OUT-X430-LSmitll_SPLITT-INt LSmitll_SPLITT

t1534 X432-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-INt 0 X432-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-IN 0 z0=5 td=1.3ps
t1535 X432-LSmitll_SPLITT-OUT-X56-LSmitll_DFFT-INt 0 X432-LSmitll_SPLITT-OUT-X56-LSmitll_DFFT-IN 0 z0=5 td=2.2ps
X432 X433-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-IN X432-LSmitll_SPLITT-OUT-X21-LSmitll_DFFT-INt X432-LSmitll_SPLITT-OUT-X56-LSmitll_DFFT-INt LSmitll_SPLITT

t1536 X433-LSmitll_SPLITT-OUT-X565-LSmitll_SPLITT-INt 0 X433-LSmitll_SPLITT-OUT-X565-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1537 X433-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-INt 0 X433-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X433 X434-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-IN X433-LSmitll_SPLITT-OUT-X565-LSmitll_SPLITT-INt X433-LSmitll_SPLITT-OUT-X432-LSmitll_SPLITT-INt LSmitll_SPLITT

t1538 X434-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-INt 0 X434-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1539 X434-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-INt 0 X434-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X434 X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-IN X434-LSmitll_SPLITT-OUT-X431-LSmitll_SPLITT-INt X434-LSmitll_SPLITT-OUT-X433-LSmitll_SPLITT-INt LSmitll_SPLITT

t1540 X435-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-INt 0 X435-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-IN 0 z0=5 td=3.2ps
t1541 X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-INt 0 X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X435 X448-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-IN X435-LSmitll_SPLITT-OUT-X429-LSmitll_SPLITT-INt X435-LSmitll_SPLITT-OUT-X434-LSmitll_SPLITT-INt LSmitll_SPLITT

t1542 X436-LSmitll_SPLITT-OUT-X66-LSmitll_AND2T-INt 0 X436-LSmitll_SPLITT-OUT-X66-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1543 X436-LSmitll_SPLITT-OUT-X305-LSmitll_OR2T-INt 0 X436-LSmitll_SPLITT-OUT-X305-LSmitll_OR2T-IN 0 z0=5 td=0.9ps
X436 X438-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-IN X436-LSmitll_SPLITT-OUT-X66-LSmitll_AND2T-INt X436-LSmitll_SPLITT-OUT-X305-LSmitll_OR2T-INt LSmitll_SPLITT

t1544 X437-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-INt 0 X437-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
t1545 X437-LSmitll_SPLITT-OUT-X282-LSmitll_AND2T-INt 0 X437-LSmitll_SPLITT-OUT-X282-LSmitll_AND2T-IN 0 z0=5 td=2.8ps
X437 X438-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-IN X437-LSmitll_SPLITT-OUT-X103-LSmitll_AND2T-INt X437-LSmitll_SPLITT-OUT-X282-LSmitll_AND2T-INt LSmitll_SPLITT

t1546 X438-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-INt 0 X438-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1547 X438-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-INt 0 X438-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X438 X441-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-IN X438-LSmitll_SPLITT-OUT-X436-LSmitll_SPLITT-INt X438-LSmitll_SPLITT-OUT-X437-LSmitll_SPLITT-INt LSmitll_SPLITT

t1548 X439-LSmitll_SPLITT-OUT-X141-LSmitll_DFFT-INt 0 X439-LSmitll_SPLITT-OUT-X141-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1549 X439-LSmitll_SPLITT-OUT-X308-LSmitll_OR2T-INt 0 X439-LSmitll_SPLITT-OUT-X308-LSmitll_OR2T-IN 0 z0=5 td=1.5ps
X439 X440-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-IN X439-LSmitll_SPLITT-OUT-X141-LSmitll_DFFT-INt X439-LSmitll_SPLITT-OUT-X308-LSmitll_OR2T-INt LSmitll_SPLITT

t1550 X440-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-INt 0 X440-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1551 X440-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-INt 0 X440-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
X440 X441-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-IN X440-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-INt X440-LSmitll_SPLITT-OUT-X439-LSmitll_SPLITT-INt LSmitll_SPLITT

t1552 X441-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-INt 0 X441-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1553 X441-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-INt 0 X441-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X441 X447-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-IN X441-LSmitll_SPLITT-OUT-X438-LSmitll_SPLITT-INt X441-LSmitll_SPLITT-OUT-X440-LSmitll_SPLITT-INt LSmitll_SPLITT

t1554 X442-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-INt 0 X442-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-IN 0 z0=5 td=0.3ps
t1555 X442-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt 0 X442-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-IN 0 z0=5 td=3.7ps
X442 X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-IN X442-LSmitll_SPLITT-OUT-X29-LSmitll_DFFT-INt X442-LSmitll_SPLITT-OUT-X104-LSmitll_AND2T-INt LSmitll_SPLITT

t1556 X443-LSmitll_SPLITT-OUT-X570-LSmitll_SPLITT-INt 0 X443-LSmitll_SPLITT-OUT-X570-LSmitll_SPLITT-IN 0 z0=5 td=1.0ps
t1557 X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-INt 0 X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X443 X446-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-IN X443-LSmitll_SPLITT-OUT-X570-LSmitll_SPLITT-INt X443-LSmitll_SPLITT-OUT-X442-LSmitll_SPLITT-INt LSmitll_SPLITT

t1558 X444-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-INt 0 X444-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1559 X444-LSmitll_SPLITT-OUT-X286-LSmitll_AND2T-INt 0 X444-LSmitll_SPLITT-OUT-X286-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
X444 X445-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-IN X444-LSmitll_SPLITT-OUT-X236-LSmitll_AND2T-INt X444-LSmitll_SPLITT-OUT-X286-LSmitll_AND2T-INt LSmitll_SPLITT

t1560 X445-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-INt 0 X445-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
t1561 X445-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-INt 0 X445-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X445 X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-IN X445-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-INt X445-LSmitll_SPLITT-OUT-X444-LSmitll_SPLITT-INt LSmitll_SPLITT

t1562 X446-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-INt 0 X446-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-IN 0 z0=5 td=5.1ps
t1563 X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-INt 0 X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X446 X447-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-IN X446-LSmitll_SPLITT-OUT-X443-LSmitll_SPLITT-INt X446-LSmitll_SPLITT-OUT-X445-LSmitll_SPLITT-INt LSmitll_SPLITT

t1564 X447-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-INt 0 X447-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1565 X447-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-INt 0 X447-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X447 X448-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-IN X447-LSmitll_SPLITT-OUT-X441-LSmitll_SPLITT-INt X447-LSmitll_SPLITT-OUT-X446-LSmitll_SPLITT-INt LSmitll_SPLITT

t1566 X448-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-INt 0 X448-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1567 X448-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-INt 0 X448-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-IN 0 z0=5 td=3.5ps
X448 X473-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-IN X448-LSmitll_SPLITT-OUT-X435-LSmitll_SPLITT-INt X448-LSmitll_SPLITT-OUT-X447-LSmitll_SPLITT-INt LSmitll_SPLITT

t1568 X449-LSmitll_SPLITT-OUT-X219-LSmitll_NDROT-INt 0 X449-LSmitll_SPLITT-OUT-X219-LSmitll_NDROT-IN 0 z0=5 td=2.6ps
t1569 X449-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-INt 0 X449-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-IN 0 z0=5 td=1.1ps
X449 X451-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-IN X449-LSmitll_SPLITT-OUT-X219-LSmitll_NDROT-INt X449-LSmitll_SPLITT-OUT-X273-LSmitll_AND2T-INt LSmitll_SPLITT

t1570 X450-LSmitll_SPLITT-OUT-X17-LSmitll_DFFT-INt 0 X450-LSmitll_SPLITT-OUT-X17-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
t1571 X450-LSmitll_SPLITT-OUT-X217-LSmitll_NDROT-INt 0 X450-LSmitll_SPLITT-OUT-X217-LSmitll_NDROT-IN 0 z0=5 td=1.7ps
X450 X451-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-IN X450-LSmitll_SPLITT-OUT-X17-LSmitll_DFFT-INt X450-LSmitll_SPLITT-OUT-X217-LSmitll_NDROT-INt LSmitll_SPLITT

t1572 X451-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-INt 0 X451-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1573 X451-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-INt 0 X451-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
X451 X454-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-IN X451-LSmitll_SPLITT-OUT-X449-LSmitll_SPLITT-INt X451-LSmitll_SPLITT-OUT-X450-LSmitll_SPLITT-INt LSmitll_SPLITT

t1574 X452-LSmitll_SPLITT-OUT-X57-LSmitll_DFFT-INt 0 X452-LSmitll_SPLITT-OUT-X57-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1575 X452-LSmitll_SPLITT-OUT-X58-LSmitll_DFFT-INt 0 X452-LSmitll_SPLITT-OUT-X58-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X452 X453-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-IN X452-LSmitll_SPLITT-OUT-X57-LSmitll_DFFT-INt X452-LSmitll_SPLITT-OUT-X58-LSmitll_DFFT-INt LSmitll_SPLITT

t1576 X453-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-INt 0 X453-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1577 X453-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-INt 0 X453-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X453 X454-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-IN X453-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-INt X453-LSmitll_SPLITT-OUT-X452-LSmitll_SPLITT-INt LSmitll_SPLITT

t1578 X454-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-INt 0 X454-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
t1579 X454-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-INt 0 X454-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X454 X460-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-IN X454-LSmitll_SPLITT-OUT-X451-LSmitll_SPLITT-INt X454-LSmitll_SPLITT-OUT-X453-LSmitll_SPLITT-INt LSmitll_SPLITT

t1580 X455-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-INt 0 X455-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1581 X455-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-INt 0 X455-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-IN 0 z0=5 td=1.9ps
X455 X456-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-IN X455-LSmitll_SPLITT-OUT-X18-LSmitll_DFFT-INt X455-LSmitll_SPLITT-OUT-X218-LSmitll_AND2T-INt LSmitll_SPLITT

t1582 X456-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-INt 0 X456-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1583 X456-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-INt 0 X456-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X456 X459-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-IN X456-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-INt X456-LSmitll_SPLITT-OUT-X455-LSmitll_SPLITT-INt LSmitll_SPLITT

t1584 X457-LSmitll_SPLITT-OUT-X53-LSmitll_DFFT-INt 0 X457-LSmitll_SPLITT-OUT-X53-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1585 X457-LSmitll_SPLITT-OUT-X54-LSmitll_DFFT-INt 0 X457-LSmitll_SPLITT-OUT-X54-LSmitll_DFFT-IN 0 z0=5 td=1.0ps
X457 X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-IN X457-LSmitll_SPLITT-OUT-X53-LSmitll_DFFT-INt X457-LSmitll_SPLITT-OUT-X54-LSmitll_DFFT-INt LSmitll_SPLITT

t1586 X458-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-INt 0 X458-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1587 X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-INt 0 X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-IN 0 z0=5 td=1.0ps
X458 X459-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-IN X458-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-INt X458-LSmitll_SPLITT-OUT-X457-LSmitll_SPLITT-INt LSmitll_SPLITT

t1588 X459-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-INt 0 X459-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-IN 0 z0=5 td=2.7ps
t1589 X459-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-INt 0 X459-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X459 X460-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-IN X459-LSmitll_SPLITT-OUT-X456-LSmitll_SPLITT-INt X459-LSmitll_SPLITT-OUT-X458-LSmitll_SPLITT-INt LSmitll_SPLITT

t1590 X460-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-INt 0 X460-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1591 X460-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-INt 0 X460-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
X460 X472-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-IN X460-LSmitll_SPLITT-OUT-X454-LSmitll_SPLITT-INt X460-LSmitll_SPLITT-OUT-X459-LSmitll_SPLITT-INt LSmitll_SPLITT

t1592 X461-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-INt 0 X461-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-IN 0 z0=5 td=6.7ps
t1593 X461-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-INt 0 X461-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-IN 0 z0=5 td=0.4ps
X461 X462-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-IN X461-LSmitll_SPLITT-OUT-X92-LSmitll_DFFT-INt X461-LSmitll_SPLITT-OUT-X281-LSmitll_AND2T-INt LSmitll_SPLITT

t1594 X462-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-INt 0 X462-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1595 X462-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-INt 0 X462-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X462 X465-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-IN X462-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-INt X462-LSmitll_SPLITT-OUT-X461-LSmitll_SPLITT-INt LSmitll_SPLITT

t1596 X463-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-INt 0 X463-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-IN 0 z0=5 td=0.2ps
t1597 X463-LSmitll_SPLITT-OUT-X237-LSmitll_NDROT-INt 0 X463-LSmitll_SPLITT-OUT-X237-LSmitll_NDROT-IN 0 z0=5 td=2.7ps
X463 X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-IN X463-LSmitll_SPLITT-OUT-X224-LSmitll_AND2T-INt X463-LSmitll_SPLITT-OUT-X237-LSmitll_NDROT-INt LSmitll_SPLITT

t1598 X464-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-INt 0 X464-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1599 X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-INt 0 X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-IN 0 z0=5 td=1.0ps
X464 X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-IN X464-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-INt X464-LSmitll_SPLITT-OUT-X463-LSmitll_SPLITT-INt LSmitll_SPLITT

t1600 X465-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-INt 0 X465-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
t1601 X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-INt 0 X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
X465 X471-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-IN X465-LSmitll_SPLITT-OUT-X462-LSmitll_SPLITT-INt X465-LSmitll_SPLITT-OUT-X464-LSmitll_SPLITT-INt LSmitll_SPLITT

t1602 X466-LSmitll_SPLITT-OUT-X93-LSmitll_DFFT-INt 0 X466-LSmitll_SPLITT-OUT-X93-LSmitll_DFFT-IN 0 z0=5 td=2.6ps
t1603 X466-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-INt 0 X466-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-IN 0 z0=5 td=1.1ps
X466 X467-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-IN X466-LSmitll_SPLITT-OUT-X93-LSmitll_DFFT-INt X466-LSmitll_SPLITT-OUT-X222-LSmitll_AND2T-INt LSmitll_SPLITT

t1604 X467-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-INt 0 X467-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-IN 0 z0=5 td=1.4ps
t1605 X467-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-INt 0 X467-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X467 X470-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-IN X467-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-INt X467-LSmitll_SPLITT-OUT-X466-LSmitll_SPLITT-INt LSmitll_SPLITT

t1606 X468-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-INt 0 X468-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1607 X468-LSmitll_SPLITT-OUT-X90-LSmitll_DFFT-INt 0 X468-LSmitll_SPLITT-OUT-X90-LSmitll_DFFT-IN 0 z0=5 td=2.0ps
X468 X469-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-IN X468-LSmitll_SPLITT-OUT-X89-LSmitll_DFFT-INt X468-LSmitll_SPLITT-OUT-X90-LSmitll_DFFT-INt LSmitll_SPLITT

t1608 X469-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-INt 0 X469-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
t1609 X469-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-INt 0 X469-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X469 X470-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-IN X469-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-INt X469-LSmitll_SPLITT-OUT-X468-LSmitll_SPLITT-INt LSmitll_SPLITT

t1610 X470-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-INt 0 X470-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
t1611 X470-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-INt 0 X470-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X470 X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-IN X470-LSmitll_SPLITT-OUT-X467-LSmitll_SPLITT-INt X470-LSmitll_SPLITT-OUT-X469-LSmitll_SPLITT-INt LSmitll_SPLITT

t1612 X471-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-INt 0 X471-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
t1613 X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-INt 0 X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X471 X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-IN X471-LSmitll_SPLITT-OUT-X465-LSmitll_SPLITT-INt X471-LSmitll_SPLITT-OUT-X470-LSmitll_SPLITT-INt LSmitll_SPLITT

t1614 X472-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-INt 0 X472-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
t1615 X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-INt 0 X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-IN 0 z0=5 td=2.8ps
X472 X473-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-IN X472-LSmitll_SPLITT-OUT-X460-LSmitll_SPLITT-INt X472-LSmitll_SPLITT-OUT-X471-LSmitll_SPLITT-INt LSmitll_SPLITT

t1616 X473-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-INt 0 X473-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-IN 0 z0=5 td=5.0ps
t1617 X473-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-INt 0 X473-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
X473 X524-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-IN X473-LSmitll_SPLITT-OUT-X448-LSmitll_SPLITT-INt X473-LSmitll_SPLITT-OUT-X472-LSmitll_SPLITT-INt LSmitll_SPLITT

t1618 X474-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-INt 0 X474-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
t1619 X474-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-INt 0 X474-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
X474 X476-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-IN X474-LSmitll_SPLITT-OUT-X140-LSmitll_DFFT-INt X474-LSmitll_SPLITT-OUT-X254-LSmitll_AND2T-INt LSmitll_SPLITT

t1620 X475-LSmitll_SPLITT-OUT-X307-LSmitll_OR2T-INt 0 X475-LSmitll_SPLITT-OUT-X307-LSmitll_OR2T-IN 0 z0=5 td=0.3ps
t1621 X475-LSmitll_SPLITT-OUT-X318-LSmitll_OR2T-INt 0 X475-LSmitll_SPLITT-OUT-X318-LSmitll_OR2T-IN 0 z0=5 td=1.5ps
X475 X476-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-IN X475-LSmitll_SPLITT-OUT-X307-LSmitll_OR2T-INt X475-LSmitll_SPLITT-OUT-X318-LSmitll_OR2T-INt LSmitll_SPLITT

t1622 X476-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-INt 0 X476-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
t1623 X476-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-INt 0 X476-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X476 X479-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-IN X476-LSmitll_SPLITT-OUT-X474-LSmitll_SPLITT-INt X476-LSmitll_SPLITT-OUT-X475-LSmitll_SPLITT-INt LSmitll_SPLITT

t1624 X477-LSmitll_SPLITT-OUT-X255-LSmitll_NDROT-INt 0 X477-LSmitll_SPLITT-OUT-X255-LSmitll_NDROT-IN 0 z0=5 td=2.2ps
t1625 X477-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-INt 0 X477-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-IN 0 z0=5 td=1.6ps
X477 X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-IN X477-LSmitll_SPLITT-OUT-X255-LSmitll_NDROT-INt X477-LSmitll_SPLITT-OUT-X256-LSmitll_AND2T-INt LSmitll_SPLITT

t1626 X478-LSmitll_SPLITT-OUT-X575-LSmitll_SPLITT-INt 0 X478-LSmitll_SPLITT-OUT-X575-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1627 X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-INt 0 X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X478 X479-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-IN X478-LSmitll_SPLITT-OUT-X575-LSmitll_SPLITT-INt X478-LSmitll_SPLITT-OUT-X477-LSmitll_SPLITT-INt LSmitll_SPLITT

t1628 X479-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-INt 0 X479-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
t1629 X479-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-INt 0 X479-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-IN 0 z0=5 td=2.2ps
X479 X485-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-IN X479-LSmitll_SPLITT-OUT-X476-LSmitll_SPLITT-INt X479-LSmitll_SPLITT-OUT-X478-LSmitll_SPLITT-INt LSmitll_SPLITT

t1630 X480-LSmitll_SPLITT-OUT-X163-LSmitll_DFFT-INt 0 X480-LSmitll_SPLITT-OUT-X163-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
t1631 X480-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-INt 0 X480-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-IN 0 z0=5 td=2.4ps
X480 X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-IN X480-LSmitll_SPLITT-OUT-X163-LSmitll_DFFT-INt X480-LSmitll_SPLITT-OUT-X285-LSmitll_AND2T-INt LSmitll_SPLITT

t1632 X481-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-INt 0 X481-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1633 X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-INt 0 X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-IN 0 z0=5 td=1.8ps
X481 X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-IN X481-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-INt X481-LSmitll_SPLITT-OUT-X480-LSmitll_SPLITT-INt LSmitll_SPLITT

t1634 X482-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-INt 0 X482-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-IN 0 z0=5 td=1.9ps
t1635 X482-LSmitll_SPLITT-OUT-X314-LSmitll_OR2T-INt 0 X482-LSmitll_SPLITT-OUT-X314-LSmitll_OR2T-IN 0 z0=5 td=3.3ps
X482 X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-IN X482-LSmitll_SPLITT-OUT-X164-LSmitll_DFFT-INt X482-LSmitll_SPLITT-OUT-X314-LSmitll_OR2T-INt LSmitll_SPLITT

t1636 X483-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-INt 0 X483-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-IN 0 z0=5 td=4.6ps
t1637 X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-INt 0 X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X483 X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-IN X483-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-INt X483-LSmitll_SPLITT-OUT-X482-LSmitll_SPLITT-INt LSmitll_SPLITT

t1638 X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-INt 0 X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1639 X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-INt 0 X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X484 X485-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-IN X484-LSmitll_SPLITT-OUT-X481-LSmitll_SPLITT-INt X484-LSmitll_SPLITT-OUT-X483-LSmitll_SPLITT-INt LSmitll_SPLITT

t1640 X485-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-INt 0 X485-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-IN 0 z0=5 td=1.5ps
t1641 X485-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-INt 0 X485-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X485 X498-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-IN X485-LSmitll_SPLITT-OUT-X479-LSmitll_SPLITT-INt X485-LSmitll_SPLITT-OUT-X484-LSmitll_SPLITT-INt LSmitll_SPLITT

t1642 X486-LSmitll_SPLITT-OUT-X295-LSmitll_AND2T-INt 0 X486-LSmitll_SPLITT-OUT-X295-LSmitll_AND2T-IN 0 z0=5 td=1.8ps
t1643 X486-LSmitll_SPLITT-OUT-X311-LSmitll_OR2T-INt 0 X486-LSmitll_SPLITT-OUT-X311-LSmitll_OR2T-IN 0 z0=5 td=1.8ps
X486 X488-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-IN X486-LSmitll_SPLITT-OUT-X295-LSmitll_AND2T-INt X486-LSmitll_SPLITT-OUT-X311-LSmitll_OR2T-INt LSmitll_SPLITT

t1644 X487-LSmitll_SPLITT-OUT-X229-LSmitll_NDROT-INt 0 X487-LSmitll_SPLITT-OUT-X229-LSmitll_NDROT-IN 0 z0=5 td=1.9ps
t1645 X487-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-INt 0 X487-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-IN 0 z0=5 td=1.2ps
X487 X488-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-IN X487-LSmitll_SPLITT-OUT-X229-LSmitll_NDROT-INt X487-LSmitll_SPLITT-OUT-X230-LSmitll_AND2T-INt LSmitll_SPLITT

t1646 X488-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-INt 0 X488-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-IN 0 z0=5 td=0.8ps
t1647 X488-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-INt 0 X488-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X488 X491-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-IN X488-LSmitll_SPLITT-OUT-X486-LSmitll_SPLITT-INt X488-LSmitll_SPLITT-OUT-X487-LSmitll_SPLITT-INt LSmitll_SPLITT

t1648 X489-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-INt 0 X489-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-IN 0 z0=5 td=3.2ps
t1649 X489-LSmitll_SPLITT-OUT-X298-LSmitll_AND2T-INt 0 X489-LSmitll_SPLITT-OUT-X298-LSmitll_AND2T-IN 0 z0=5 td=3.9ps
X489 X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-IN X489-LSmitll_SPLITT-OUT-X35-LSmitll_OR2T-INt X489-LSmitll_SPLITT-OUT-X298-LSmitll_AND2T-INt LSmitll_SPLITT

t1650 X490-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-INt 0 X490-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
t1651 X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-INt 0 X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X490 X491-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-IN X490-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-INt X490-LSmitll_SPLITT-OUT-X489-LSmitll_SPLITT-INt LSmitll_SPLITT

t1652 X491-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-INt 0 X491-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-IN 0 z0=5 td=0.5ps
t1653 X491-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-INt 0 X491-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
X491 X497-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-IN X491-LSmitll_SPLITT-OUT-X488-LSmitll_SPLITT-INt X491-LSmitll_SPLITT-OUT-X490-LSmitll_SPLITT-INt LSmitll_SPLITT

t1654 X492-LSmitll_SPLITT-OUT-X294-LSmitll_AND2T-INt 0 X492-LSmitll_SPLITT-OUT-X294-LSmitll_AND2T-IN 0 z0=5 td=7.4ps
t1655 X492-LSmitll_SPLITT-OUT-X321-LSmitll_OR2T-INt 0 X492-LSmitll_SPLITT-OUT-X321-LSmitll_OR2T-IN 0 z0=5 td=2.9ps
X492 X493-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-IN X492-LSmitll_SPLITT-OUT-X294-LSmitll_AND2T-INt X492-LSmitll_SPLITT-OUT-X321-LSmitll_OR2T-INt LSmitll_SPLITT

t1656 X493-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-INt 0 X493-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1657 X493-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-INt 0 X493-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X493 X496-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-IN X493-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-INt X493-LSmitll_SPLITT-OUT-X492-LSmitll_SPLITT-INt LSmitll_SPLITT

t1658 X494-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-INt 0 X494-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-IN 0 z0=5 td=3.1ps
t1659 X494-LSmitll_SPLITT-OUT-X244-LSmitll_AND2T-INt 0 X494-LSmitll_SPLITT-OUT-X244-LSmitll_AND2T-IN 0 z0=5 td=3.0ps
X494 X495-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-IN X494-LSmitll_SPLITT-OUT-X36-LSmitll_OR2T-INt X494-LSmitll_SPLITT-OUT-X244-LSmitll_AND2T-INt LSmitll_SPLITT

t1660 X495-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-INt 0 X495-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
t1661 X495-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-INt 0 X495-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X495 X496-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-IN X495-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-INt X495-LSmitll_SPLITT-OUT-X494-LSmitll_SPLITT-INt LSmitll_SPLITT

t1662 X496-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-INt 0 X496-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1663 X496-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-INt 0 X496-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
X496 X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-IN X496-LSmitll_SPLITT-OUT-X493-LSmitll_SPLITT-INt X496-LSmitll_SPLITT-OUT-X495-LSmitll_SPLITT-INt LSmitll_SPLITT

t1664 X497-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-INt 0 X497-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1665 X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-INt 0 X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-IN 0 z0=5 td=1.3ps
X497 X498-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-IN X497-LSmitll_SPLITT-OUT-X491-LSmitll_SPLITT-INt X497-LSmitll_SPLITT-OUT-X496-LSmitll_SPLITT-INt LSmitll_SPLITT

t1666 X498-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-INt 0 X498-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-IN 0 z0=5 td=4.1ps
t1667 X498-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-INt 0 X498-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X498 X523-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-IN X498-LSmitll_SPLITT-OUT-X485-LSmitll_SPLITT-INt X498-LSmitll_SPLITT-OUT-X497-LSmitll_SPLITT-INt LSmitll_SPLITT

t1668 X499-LSmitll_SPLITT-OUT-X225-LSmitll_NDROT-INt 0 X499-LSmitll_SPLITT-OUT-X225-LSmitll_NDROT-IN 0 z0=5 td=2.2ps
t1669 X499-LSmitll_SPLITT-OUT-X289-LSmitll_AND2T-INt 0 X499-LSmitll_SPLITT-OUT-X289-LSmitll_AND2T-IN 0 z0=5 td=0.4ps
X499 X501-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-IN X499-LSmitll_SPLITT-OUT-X225-LSmitll_NDROT-INt X499-LSmitll_SPLITT-OUT-X289-LSmitll_AND2T-INt LSmitll_SPLITT

t1670 X500-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-INt 0 X500-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-IN 0 z0=5 td=0.4ps
t1671 X500-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-INt 0 X500-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-IN 0 z0=5 td=2.5ps
X500 X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-IN X500-LSmitll_SPLITT-OUT-X183-LSmitll_DFFT-INt X500-LSmitll_SPLITT-OUT-X226-LSmitll_AND2T-INt LSmitll_SPLITT

t1672 X501-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-INt 0 X501-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1673 X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-INt 0 X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-IN 0 z0=5 td=1.7ps
X501 X504-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-IN X501-LSmitll_SPLITT-OUT-X499-LSmitll_SPLITT-INt X501-LSmitll_SPLITT-OUT-X500-LSmitll_SPLITT-INt LSmitll_SPLITT

t1674 X502-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-INt 0 X502-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-IN 0 z0=5 td=3.1ps
t1675 X502-LSmitll_SPLITT-OUT-X299-LSmitll_AND2T-INt 0 X502-LSmitll_SPLITT-OUT-X299-LSmitll_AND2T-IN 0 z0=5 td=1.3ps
X502 X503-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-IN X502-LSmitll_SPLITT-OUT-X184-LSmitll_DFFT-INt X502-LSmitll_SPLITT-OUT-X299-LSmitll_AND2T-INt LSmitll_SPLITT

t1676 X503-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-INt 0 X503-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-IN 0 z0=5 td=3.0ps
t1677 X503-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-INt 0 X503-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-IN 0 z0=5 td=1.9ps
X503 X504-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-IN X503-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-INt X503-LSmitll_SPLITT-OUT-X502-LSmitll_SPLITT-INt LSmitll_SPLITT

t1678 X504-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-INt 0 X504-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-IN 0 z0=5 td=0.5ps
t1679 X504-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-INt 0 X504-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
X504 X510-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-IN X504-LSmitll_SPLITT-OUT-X501-LSmitll_SPLITT-INt X504-LSmitll_SPLITT-OUT-X503-LSmitll_SPLITT-INt LSmitll_SPLITT

t1680 X505-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-INt 0 X505-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-IN 0 z0=5 td=4.7ps
t1681 X505-LSmitll_SPLITT-OUT-X185-LSmitll_DFFT-INt 0 X505-LSmitll_SPLITT-OUT-X185-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
X505 X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-IN X505-LSmitll_SPLITT-OUT-X138-LSmitll_DFFT-INt X505-LSmitll_SPLITT-OUT-X185-LSmitll_DFFT-INt LSmitll_SPLITT

t1682 X506-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-INt 0 X506-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
t1683 X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-INt 0 X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
X506 X509-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-IN X506-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-INt X506-LSmitll_SPLITT-OUT-X505-LSmitll_SPLITT-INt LSmitll_SPLITT

t1684 X507-LSmitll_SPLITT-OUT-X157-LSmitll_DFFT-INt 0 X507-LSmitll_SPLITT-OUT-X157-LSmitll_DFFT-IN 0 z0=5 td=2.0ps
t1685 X507-LSmitll_SPLITT-OUT-X158-LSmitll_DFFT-INt 0 X507-LSmitll_SPLITT-OUT-X158-LSmitll_DFFT-IN 0 z0=5 td=3.2ps
X507 X508-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-IN X507-LSmitll_SPLITT-OUT-X157-LSmitll_DFFT-INt X507-LSmitll_SPLITT-OUT-X158-LSmitll_DFFT-INt LSmitll_SPLITT

t1686 X508-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-INt 0 X508-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1687 X508-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-INt 0 X508-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-IN 0 z0=5 td=2.9ps
X508 X509-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-IN X508-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-INt X508-LSmitll_SPLITT-OUT-X507-LSmitll_SPLITT-INt LSmitll_SPLITT

t1688 X509-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-INt 0 X509-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-IN 0 z0=5 td=0.9ps
t1689 X509-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-INt 0 X509-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-IN 0 z0=5 td=0.7ps
X509 X510-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-IN X509-LSmitll_SPLITT-OUT-X506-LSmitll_SPLITT-INt X509-LSmitll_SPLITT-OUT-X508-LSmitll_SPLITT-INt LSmitll_SPLITT

t1690 X510-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-INt 0 X510-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-IN 0 z0=5 td=3.3ps
t1691 X510-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-INt 0 X510-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
X510 X522-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-IN X510-LSmitll_SPLITT-OUT-X504-LSmitll_SPLITT-INt X510-LSmitll_SPLITT-OUT-X509-LSmitll_SPLITT-INt LSmitll_SPLITT

t1692 X511-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-INt 0 X511-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-IN 0 z0=5 td=0.9ps
t1693 X511-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-INt 0 X511-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-IN 0 z0=5 td=1.1ps
X511 X512-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-IN X511-LSmitll_SPLITT-OUT-X177-LSmitll_DFFT-INt X511-LSmitll_SPLITT-OUT-X178-LSmitll_DFFT-INt LSmitll_SPLITT

t1694 X512-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-INt 0 X512-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-IN 0 z0=5 td=2.4ps
t1695 X512-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-INt 0 X512-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
X512 X515-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-IN X512-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-INt X512-LSmitll_SPLITT-OUT-X511-LSmitll_SPLITT-INt LSmitll_SPLITT

t1696 X513-LSmitll_SPLITT-OUT-X72-LSmitll_AND2T-INt 0 X513-LSmitll_SPLITT-OUT-X72-LSmitll_AND2T-IN 0 z0=5 td=0.7ps
t1697 X513-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-INt 0 X513-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-IN 0 z0=5 td=2.3ps
X513 X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-IN X513-LSmitll_SPLITT-OUT-X72-LSmitll_AND2T-INt X513-LSmitll_SPLITT-OUT-X160-LSmitll_DFFT-INt LSmitll_SPLITT

t1698 X514-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-INt 0 X514-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-IN 0 z0=5 td=1.0ps
t1699 X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-INt 0 X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-IN 0 z0=5 td=1.0ps
X514 X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-IN X514-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-INt X514-LSmitll_SPLITT-OUT-X513-LSmitll_SPLITT-INt LSmitll_SPLITT

t1700 X515-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-INt 0 X515-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
t1701 X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-INt 0 X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-IN 0 z0=5 td=2.1ps
X515 X521-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-IN X515-LSmitll_SPLITT-OUT-X512-LSmitll_SPLITT-INt X515-LSmitll_SPLITT-OUT-X514-LSmitll_SPLITT-INt LSmitll_SPLITT

t1702 X516-LSmitll_SPLITT-OUT-X227-LSmitll_NDROT-INt 0 X516-LSmitll_SPLITT-OUT-X227-LSmitll_NDROT-IN 0 z0=5 td=1.9ps
t1703 X516-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-INt 0 X516-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-IN 0 z0=5 td=2.7ps
X516 X517-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-IN X516-LSmitll_SPLITT-OUT-X227-LSmitll_NDROT-INt X516-LSmitll_SPLITT-OUT-X242-LSmitll_AND2T-INt LSmitll_SPLITT

t1704 X517-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-INt 0 X517-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1705 X517-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-INt 0 X517-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-IN 0 z0=5 td=1.1ps
X517 X520-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-IN X517-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-INt X517-LSmitll_SPLITT-OUT-X516-LSmitll_SPLITT-INt LSmitll_SPLITT

t1706 X518-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-INt 0 X518-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-IN 0 z0=5 td=1.6ps
t1707 X518-LSmitll_SPLITT-OUT-X241-LSmitll_NDROT-INt 0 X518-LSmitll_SPLITT-OUT-X241-LSmitll_NDROT-IN 0 z0=5 td=2.0ps
X518 X519-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-IN X518-LSmitll_SPLITT-OUT-X32-LSmitll_DFFT-INt X518-LSmitll_SPLITT-OUT-X241-LSmitll_NDROT-INt LSmitll_SPLITT

t1708 X519-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-INt 0 X519-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-IN 0 z0=5 td=2.0ps
t1709 X519-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-INt 0 X519-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-IN 0 z0=5 td=2.5ps
X519 X520-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-IN X519-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-INt X519-LSmitll_SPLITT-OUT-X518-LSmitll_SPLITT-INt LSmitll_SPLITT

t1710 X520-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-INt 0 X520-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-IN 0 z0=5 td=3.5ps
t1711 X520-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-INt 0 X520-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-IN 0 z0=5 td=2.3ps
X520 X521-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-IN X520-LSmitll_SPLITT-OUT-X517-LSmitll_SPLITT-INt X520-LSmitll_SPLITT-OUT-X519-LSmitll_SPLITT-INt LSmitll_SPLITT

t1712 X521-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-INt 0 X521-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-IN 0 z0=5 td=1.6ps
t1713 X521-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-INt 0 X521-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-IN 0 z0=5 td=1.2ps
X521 X522-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-IN X521-LSmitll_SPLITT-OUT-X515-LSmitll_SPLITT-INt X521-LSmitll_SPLITT-OUT-X520-LSmitll_SPLITT-INt LSmitll_SPLITT

t1714 X522-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-INt 0 X522-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-IN 0 z0=5 td=3.1ps
t1715 X522-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-INt 0 X522-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-IN 0 z0=5 td=3.4ps
X522 X523-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-IN X522-LSmitll_SPLITT-OUT-X510-LSmitll_SPLITT-INt X522-LSmitll_SPLITT-OUT-X521-LSmitll_SPLITT-INt LSmitll_SPLITT

t1716 X523-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-INt 0 X523-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-IN 0 z0=5 td=3.8ps
t1717 X523-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-INt 0 X523-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-IN 0 z0=5 td=4.6ps
X523 X524-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-IN X523-LSmitll_SPLITT-OUT-X498-LSmitll_SPLITT-INt X523-LSmitll_SPLITT-OUT-X522-LSmitll_SPLITT-INt LSmitll_SPLITT

t1718 X524-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-INt 0 X524-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-IN 0 z0=5 td=6.5ps
t1719 X524-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-INt 0 X524-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-IN 0 z0=5 td=4.7ps
X524 X576-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-IN X524-LSmitll_SPLITT-OUT-X473-LSmitll_SPLITT-INt X524-LSmitll_SPLITT-OUT-X523-LSmitll_SPLITT-INt LSmitll_SPLITT

t1720 X525-LSmitll_SPLITT-OUT-X19-LSmitll_DFFT-INt 0 X525-LSmitll_SPLITT-OUT-X19-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1721 X525-SPLITT-OUT-R-INt 0 X525-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X525 X456-LSmitll_SPLITT-OUT-X525-LSmitll_SPLITT-IN X525-LSmitll_SPLITT-OUT-X19-LSmitll_DFFT-INt X525-SPLITT-OUT-R-INt LSmitll_SPLITT

t1722 X526-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-INt 0 X526-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-IN 0 z0=5 td=1.2ps
t1723 X526-SPLITT-OUT-R-INt 0 X526-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X526 X418-LSmitll_SPLITT-OUT-X526-LSmitll_SPLITT-IN X526-LSmitll_SPLITT-OUT-X33-LSmitll_OR2T-INt X526-SPLITT-OUT-R-INt LSmitll_SPLITT

t1724 X527-LSmitll_SPLITT-OUT-X38-LSmitll_NOTT-INt 0 X527-LSmitll_SPLITT-OUT-X38-LSmitll_NOTT-IN 0 z0=5 td=0.3ps
t1725 X527-SPLITT-OUT-R-INt 0 X527-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X527 X338-LSmitll_SPLITT-OUT-X527-LSmitll_SPLITT-IN X527-LSmitll_SPLITT-OUT-X38-LSmitll_NOTT-INt X527-SPLITT-OUT-R-INt LSmitll_SPLITT

t1726 X528-LSmitll_SPLITT-OUT-X40-LSmitll_NOTT-INt 0 X528-LSmitll_SPLITT-OUT-X40-LSmitll_NOTT-IN 0 z0=5 td=0.9ps
t1727 X528-SPLITT-OUT-R-INt 0 X528-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X528 X519-LSmitll_SPLITT-OUT-X528-LSmitll_SPLITT-IN X528-LSmitll_SPLITT-OUT-X40-LSmitll_NOTT-INt X528-SPLITT-OUT-R-INt LSmitll_SPLITT

t1728 X529-LSmitll_SPLITT-OUT-X55-LSmitll_DFFT-INt 0 X529-LSmitll_SPLITT-OUT-X55-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1729 X529-SPLITT-OUT-R-INt 0 X529-SPLITT-OUT-R-IN 0 z0=5 td=9.9ps
X529 X458-LSmitll_SPLITT-OUT-X529-LSmitll_SPLITT-IN X529-LSmitll_SPLITT-OUT-X55-LSmitll_DFFT-INt X529-SPLITT-OUT-R-INt LSmitll_SPLITT

t1730 X530-LSmitll_SPLITT-OUT-X68-LSmitll_AND2T-INt 0 X530-LSmitll_SPLITT-OUT-X68-LSmitll_AND2T-IN 0 z0=5 td=0.5ps
t1731 X530-SPLITT-OUT-R-INt 0 X530-SPLITT-OUT-R-IN 0 z0=5 td=10.0ps
X530 X380-LSmitll_SPLITT-OUT-X530-LSmitll_SPLITT-IN X530-LSmitll_SPLITT-OUT-X68-LSmitll_AND2T-INt X530-SPLITT-OUT-R-INt LSmitll_SPLITT

t1732 X531-LSmitll_SPLITT-OUT-X69-LSmitll_AND2T-INt 0 X531-LSmitll_SPLITT-OUT-X69-LSmitll_AND2T-IN 0 z0=5 td=2.1ps
t1733 X531-SPLITT-OUT-R-INt 0 X531-SPLITT-OUT-R-IN 0 z0=5 td=9.7ps
X531 X394-LSmitll_SPLITT-OUT-X531-LSmitll_SPLITT-IN X531-LSmitll_SPLITT-OUT-X69-LSmitll_AND2T-INt X531-SPLITT-OUT-R-INt LSmitll_SPLITT

t1734 X532-LSmitll_SPLITT-OUT-X71-LSmitll_AND2T-INt 0 X532-LSmitll_SPLITT-OUT-X71-LSmitll_AND2T-IN 0 z0=5 td=0.9ps
t1735 X532-SPLITT-OUT-R-INt 0 X532-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X532 X514-LSmitll_SPLITT-OUT-X532-LSmitll_SPLITT-IN X532-LSmitll_SPLITT-OUT-X71-LSmitll_AND2T-INt X532-SPLITT-OUT-R-INt LSmitll_SPLITT

t1736 X533-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-INt 0 X533-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1737 X533-SPLITT-OUT-R-INt 0 X533-SPLITT-OUT-R-IN 0 z0=5 td=9.9ps
X533 X469-LSmitll_SPLITT-OUT-X533-LSmitll_SPLITT-IN X533-LSmitll_SPLITT-OUT-X91-LSmitll_DFFT-INt X533-SPLITT-OUT-R-INt LSmitll_SPLITT

t1738 X534-LSmitll_SPLITT-OUT-X94-LSmitll_DFFT-INt 0 X534-LSmitll_SPLITT-OUT-X94-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
t1739 X534-SPLITT-OUT-R-INt 0 X534-SPLITT-OUT-R-IN 0 z0=5 td=10.0ps
X534 X467-LSmitll_SPLITT-OUT-X534-LSmitll_SPLITT-IN X534-LSmitll_SPLITT-OUT-X94-LSmitll_DFFT-INt X534-SPLITT-OUT-R-INt LSmitll_SPLITT

t1740 X535-LSmitll_SPLITT-OUT-X97-LSmitll_DFFT-INt 0 X535-LSmitll_SPLITT-OUT-X97-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1741 X535-SPLITT-OUT-R-INt 0 X535-SPLITT-OUT-R-IN 0 z0=5 td=10.1ps
X535 X363-LSmitll_SPLITT-OUT-X535-LSmitll_SPLITT-IN X535-LSmitll_SPLITT-OUT-X97-LSmitll_DFFT-INt X535-SPLITT-OUT-R-INt LSmitll_SPLITT

t1742 X536-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-INt 0 X536-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-IN 0 z0=5 td=0.8ps
t1743 X536-SPLITT-OUT-R-INt 0 X536-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X536 X389-LSmitll_SPLITT-OUT-X536-LSmitll_SPLITT-IN X536-LSmitll_SPLITT-OUT-X105-LSmitll_AND2T-INt X536-SPLITT-OUT-R-INt LSmitll_SPLITT

t1744 X537-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-INt 0 X537-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-IN 0 z0=5 td=0.8ps
t1745 X537-SPLITT-OUT-R-INt 0 X537-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X537 X413-LSmitll_SPLITT-OUT-X537-LSmitll_SPLITT-IN X537-LSmitll_SPLITT-OUT-X106-LSmitll_AND2T-INt X537-SPLITT-OUT-R-INt LSmitll_SPLITT

t1746 X538-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt 0 X538-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-IN 0 z0=5 td=2.0ps
t1747 X538-SPLITT-OUT-R-INt 0 X538-SPLITT-OUT-R-IN 0 z0=5 td=9.8ps
X538 X392-LSmitll_SPLITT-OUT-X538-LSmitll_SPLITT-IN X538-LSmitll_SPLITT-OUT-X107-LSmitll_AND2T-INt X538-SPLITT-OUT-R-INt LSmitll_SPLITT

t1748 X539-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-INt 0 X539-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
t1749 X539-SPLITT-OUT-R-INt 0 X539-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X539 X464-LSmitll_SPLITT-OUT-X539-LSmitll_SPLITT-IN X539-LSmitll_SPLITT-OUT-X137-LSmitll_DFFT-INt X539-SPLITT-OUT-R-INt LSmitll_SPLITT

t1750 X540-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-INt 0 X540-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1751 X540-SPLITT-OUT-R-INt 0 X540-SPLITT-OUT-R-IN 0 z0=5 td=10.5ps
X540 X506-LSmitll_SPLITT-OUT-X540-LSmitll_SPLITT-IN X540-LSmitll_SPLITT-OUT-X139-LSmitll_DFFT-INt X540-SPLITT-OUT-R-INt LSmitll_SPLITT

t1752 X541-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-INt 0 X541-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
t1753 X541-SPLITT-OUT-R-INt 0 X541-SPLITT-OUT-R-IN 0 z0=5 td=9.8ps
X541 X405-LSmitll_SPLITT-OUT-X541-LSmitll_SPLITT-IN X541-LSmitll_SPLITT-OUT-X142-LSmitll_DFFT-INt X541-SPLITT-OUT-R-INt LSmitll_SPLITT

t1754 X542-LSmitll_SPLITT-OUT-X159-LSmitll_DFFT-INt 0 X542-LSmitll_SPLITT-OUT-X159-LSmitll_DFFT-IN 0 z0=5 td=0.5ps
t1755 X542-SPLITT-OUT-R-INt 0 X542-SPLITT-OUT-R-IN 0 z0=5 td=10.1ps
X542 X508-LSmitll_SPLITT-OUT-X542-LSmitll_SPLITT-IN X542-LSmitll_SPLITT-OUT-X159-LSmitll_DFFT-INt X542-SPLITT-OUT-R-INt LSmitll_SPLITT

t1756 X543-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-INt 0 X543-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1757 X543-SPLITT-OUT-R-INt 0 X543-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X543 X483-LSmitll_SPLITT-OUT-X543-LSmitll_SPLITT-IN X543-LSmitll_SPLITT-OUT-X165-LSmitll_DFFT-INt X543-SPLITT-OUT-R-INt LSmitll_SPLITT

t1758 X544-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-INt 0 X544-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-IN 0 z0=5 td=0.6ps
t1759 X544-SPLITT-OUT-R-INt 0 X544-SPLITT-OUT-R-IN 0 z0=5 td=9.5ps
X544 X382-LSmitll_SPLITT-OUT-X544-LSmitll_SPLITT-IN X544-LSmitll_SPLITT-OUT-X166-LSmitll_DFFT-INt X544-SPLITT-OUT-R-INt LSmitll_SPLITT

t1760 X545-LSmitll_SPLITT-OUT-X179-LSmitll_DFFT-INt 0 X545-LSmitll_SPLITT-OUT-X179-LSmitll_DFFT-IN 0 z0=5 td=0.7ps
t1761 X545-SPLITT-OUT-R-INt 0 X545-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X545 X493-LSmitll_SPLITT-OUT-X545-LSmitll_SPLITT-IN X545-LSmitll_SPLITT-OUT-X179-LSmitll_DFFT-INt X545-SPLITT-OUT-R-INt LSmitll_SPLITT

t1762 X546-LSmitll_SPLITT-OUT-X180-LSmitll_DFFT-INt 0 X546-LSmitll_SPLITT-OUT-X180-LSmitll_DFFT-IN 0 z0=5 td=0.8ps
t1763 X546-SPLITT-OUT-R-INt 0 X546-SPLITT-OUT-R-IN 0 z0=5 td=9.5ps
X546 X495-LSmitll_SPLITT-OUT-X546-LSmitll_SPLITT-IN X546-LSmitll_SPLITT-OUT-X180-LSmitll_DFFT-INt X546-SPLITT-OUT-R-INt LSmitll_SPLITT

t1764 X547-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-INt 0 X547-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
t1765 X547-SPLITT-OUT-R-INt 0 X547-SPLITT-OUT-R-IN 0 z0=5 td=9.8ps
X547 X453-LSmitll_SPLITT-OUT-X547-LSmitll_SPLITT-IN X547-LSmitll_SPLITT-OUT-X220-LSmitll_AND2T-INt X547-SPLITT-OUT-R-INt LSmitll_SPLITT

t1766 X548-LSmitll_SPLITT-OUT-X221-LSmitll_NDROT-INt 0 X548-LSmitll_SPLITT-OUT-X221-LSmitll_NDROT-IN 0 z0=5 td=0.9ps
t1767 X548-SPLITT-OUT-R-INt 0 X548-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X548 X462-LSmitll_SPLITT-OUT-X548-LSmitll_SPLITT-IN X548-LSmitll_SPLITT-OUT-X221-LSmitll_NDROT-INt X548-SPLITT-OUT-R-INt LSmitll_SPLITT

t1768 X549-LSmitll_SPLITT-OUT-X223-LSmitll_NDROT-INt 0 X549-LSmitll_SPLITT-OUT-X223-LSmitll_NDROT-IN 0 z0=5 td=0.8ps
t1769 X549-SPLITT-OUT-R-INt 0 X549-SPLITT-OUT-R-IN 0 z0=5 td=9.9ps
X549 X481-LSmitll_SPLITT-OUT-X549-LSmitll_SPLITT-IN X549-LSmitll_SPLITT-OUT-X223-LSmitll_NDROT-INt X549-SPLITT-OUT-R-INt LSmitll_SPLITT

t1770 X550-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-INt 0 X550-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-IN 0 z0=5 td=0.7ps
t1771 X550-SPLITT-OUT-R-INt 0 X550-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X550 X517-LSmitll_SPLITT-OUT-X550-LSmitll_SPLITT-IN X550-LSmitll_SPLITT-OUT-X228-LSmitll_AND2T-INt X550-SPLITT-OUT-R-INt LSmitll_SPLITT

t1772 X551-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-INt 0 X551-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
t1773 X551-SPLITT-OUT-R-INt 0 X551-SPLITT-OUT-R-IN 0 z0=5 td=9.7ps
X551 X431-LSmitll_SPLITT-OUT-X551-LSmitll_SPLITT-IN X551-LSmitll_SPLITT-OUT-X232-LSmitll_AND2T-INt X551-SPLITT-OUT-R-INt LSmitll_SPLITT

t1774 X552-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt 0 X552-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
t1775 X552-SPLITT-OUT-R-INt 0 X552-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X552 X428-LSmitll_SPLITT-OUT-X552-LSmitll_SPLITT-IN X552-LSmitll_SPLITT-OUT-X234-LSmitll_AND2T-INt X552-SPLITT-OUT-R-INt LSmitll_SPLITT

t1776 X553-LSmitll_SPLITT-OUT-X235-LSmitll_NDROT-INt 0 X553-LSmitll_SPLITT-OUT-X235-LSmitll_NDROT-IN 0 z0=5 td=0.7ps
t1777 X553-SPLITT-OUT-R-INt 0 X553-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X553 X440-LSmitll_SPLITT-OUT-X553-LSmitll_SPLITT-IN X553-LSmitll_SPLITT-OUT-X235-LSmitll_NDROT-INt X553-SPLITT-OUT-R-INt LSmitll_SPLITT

t1778 X554-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt 0 X554-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
t1779 X554-SPLITT-OUT-R-INt 0 X554-SPLITT-OUT-R-IN 0 z0=5 td=10.2ps
X554 X445-LSmitll_SPLITT-OUT-X554-LSmitll_SPLITT-IN X554-LSmitll_SPLITT-OUT-X238-LSmitll_AND2T-INt X554-SPLITT-OUT-R-INt LSmitll_SPLITT

t1780 X555-LSmitll_SPLITT-OUT-X243-LSmitll_NDROT-INt 0 X555-LSmitll_SPLITT-OUT-X243-LSmitll_NDROT-IN 0 z0=5 td=1.3ps
t1781 X555-SPLITT-OUT-R-INt 0 X555-SPLITT-OUT-R-IN 0 z0=5 td=9.8ps
X555 X490-LSmitll_SPLITT-OUT-X555-LSmitll_SPLITT-IN X555-LSmitll_SPLITT-OUT-X243-LSmitll_NDROT-INt X555-SPLITT-OUT-R-INt LSmitll_SPLITT

t1782 X556-LSmitll_SPLITT-OUT-X245-LSmitll_NDROT-INt 0 X556-LSmitll_SPLITT-OUT-X245-LSmitll_NDROT-IN 0 z0=5 td=0.9ps
t1783 X556-SPLITT-OUT-R-INt 0 X556-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X556 X354-LSmitll_SPLITT-OUT-X556-LSmitll_SPLITT-IN X556-LSmitll_SPLITT-OUT-X245-LSmitll_NDROT-INt X556-SPLITT-OUT-R-INt LSmitll_SPLITT

t1784 X557-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-INt 0 X557-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
t1785 X557-SPLITT-OUT-R-INt 0 X557-SPLITT-OUT-R-IN 0 z0=5 td=9.8ps
X557 X366-LSmitll_SPLITT-OUT-X557-LSmitll_SPLITT-IN X557-LSmitll_SPLITT-OUT-X250-LSmitll_AND2T-INt X557-SPLITT-OUT-R-INt LSmitll_SPLITT

t1786 X558-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-INt 0 X558-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
t1787 X558-SPLITT-OUT-R-INt 0 X558-SPLITT-OUT-R-IN 0 z0=5 td=10.1ps
X558 X368-LSmitll_SPLITT-OUT-X558-LSmitll_SPLITT-IN X558-LSmitll_SPLITT-OUT-X252-LSmitll_AND2T-INt X558-SPLITT-OUT-R-INt LSmitll_SPLITT

t1788 X559-LSmitll_SPLITT-OUT-X253-LSmitll_NDROT-INt 0 X559-LSmitll_SPLITT-OUT-X253-LSmitll_NDROT-IN 0 z0=5 td=0.9ps
t1789 X559-SPLITT-OUT-R-INt 0 X559-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X559 X407-LSmitll_SPLITT-OUT-X559-LSmitll_SPLITT-IN X559-LSmitll_SPLITT-OUT-X253-LSmitll_NDROT-INt X559-SPLITT-OUT-R-INt LSmitll_SPLITT

t1790 X560-LSmitll_SPLITT-OUT-X257-LSmitll_NDROT-INt 0 X560-LSmitll_SPLITT-OUT-X257-LSmitll_NDROT-IN 0 z0=5 td=1.0ps
t1791 X560-SPLITT-OUT-R-INt 0 X560-SPLITT-OUT-R-IN 0 z0=5 td=10.1ps
X560 X512-LSmitll_SPLITT-OUT-X560-LSmitll_SPLITT-IN X560-LSmitll_SPLITT-OUT-X257-LSmitll_NDROT-INt X560-SPLITT-OUT-R-INt LSmitll_SPLITT

t1792 X561-LSmitll_SPLITT-OUT-X258-LSmitll_AND2T-INt 0 X561-LSmitll_SPLITT-OUT-X258-LSmitll_AND2T-IN 0 z0=5 td=1.0ps
t1793 X561-SPLITT-OUT-R-INt 0 X561-SPLITT-OUT-R-IN 0 z0=5 td=9.9ps
X561 X503-LSmitll_SPLITT-OUT-X561-LSmitll_SPLITT-IN X561-LSmitll_SPLITT-OUT-X258-LSmitll_AND2T-INt X561-SPLITT-OUT-R-INt LSmitll_SPLITT

t1794 X562-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-INt 0 X562-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
t1795 X562-SPLITT-OUT-R-INt 0 X562-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X562 X329-LSmitll_SPLITT-OUT-X562-LSmitll_SPLITT-IN X562-LSmitll_SPLITT-OUT-X260-LSmitll_AND2T-INt X562-SPLITT-OUT-R-INt LSmitll_SPLITT

t1796 X563-LSmitll_SPLITT-OUT-X263-LSmitll_NDROT-INt 0 X563-LSmitll_SPLITT-OUT-X263-LSmitll_NDROT-IN 0 z0=5 td=0.9ps
t1797 X563-SPLITT-OUT-R-INt 0 X563-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X563 X341-LSmitll_SPLITT-OUT-X563-LSmitll_SPLITT-IN X563-LSmitll_SPLITT-OUT-X263-LSmitll_NDROT-INt X563-SPLITT-OUT-R-INt LSmitll_SPLITT

t1798 X564-LSmitll_SPLITT-OUT-X271-LSmitll_NDROT-INt 0 X564-LSmitll_SPLITT-OUT-X271-LSmitll_NDROT-IN 0 z0=5 td=1.2ps
t1799 X564-SPLITT-OUT-R-INt 0 X564-SPLITT-OUT-R-IN 0 z0=5 td=10.1ps
X564 X377-LSmitll_SPLITT-OUT-X564-LSmitll_SPLITT-IN X564-LSmitll_SPLITT-OUT-X271-LSmitll_NDROT-INt X564-SPLITT-OUT-R-INt LSmitll_SPLITT

t1800 X565-LSmitll_SPLITT-OUT-X277-LSmitll_AND2T-INt 0 X565-LSmitll_SPLITT-OUT-X277-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
t1801 X565-SPLITT-OUT-R-INt 0 X565-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X565 X433-LSmitll_SPLITT-OUT-X565-LSmitll_SPLITT-IN X565-LSmitll_SPLITT-OUT-X277-LSmitll_AND2T-INt X565-SPLITT-OUT-R-INt LSmitll_SPLITT

t1802 X566-LSmitll_SPLITT-OUT-X280-LSmitll_AND2T-INt 0 X566-LSmitll_SPLITT-OUT-X280-LSmitll_AND2T-IN 0 z0=5 td=0.6ps
t1803 X566-SPLITT-OUT-R-INt 0 X566-SPLITT-OUT-R-IN 0 z0=5 td=10.1ps
X566 X326-LSmitll_SPLITT-OUT-X566-LSmitll_SPLITT-IN X566-LSmitll_SPLITT-OUT-X280-LSmitll_AND2T-INt X566-SPLITT-OUT-R-INt LSmitll_SPLITT

t1804 X567-LSmitll_SPLITT-OUT-X283-LSmitll_AND2T-INt 0 X567-LSmitll_SPLITT-OUT-X283-LSmitll_AND2T-IN 0 z0=5 td=0.4ps
t1805 X567-SPLITT-OUT-R-INt 0 X567-SPLITT-OUT-R-IN 0 z0=5 td=9.5ps
X567 X331-LSmitll_SPLITT-OUT-X567-LSmitll_SPLITT-IN X567-LSmitll_SPLITT-OUT-X283-LSmitll_AND2T-INt X567-SPLITT-OUT-R-INt LSmitll_SPLITT

t1806 X568-LSmitll_SPLITT-OUT-X297-LSmitll_AND2T-INt 0 X568-LSmitll_SPLITT-OUT-X297-LSmitll_AND2T-IN 0 z0=5 td=0.5ps
t1807 X568-SPLITT-OUT-R-INt 0 X568-SPLITT-OUT-R-IN 0 z0=5 td=10.4ps
X568 X411-LSmitll_SPLITT-OUT-X568-LSmitll_SPLITT-IN X568-LSmitll_SPLITT-OUT-X297-LSmitll_AND2T-INt X568-SPLITT-OUT-R-INt LSmitll_SPLITT

t1808 X569-LSmitll_SPLITT-OUT-X301-LSmitll_OR2T-INt 0 X569-LSmitll_SPLITT-OUT-X301-LSmitll_OR2T-IN 0 z0=5 td=0.7ps
t1809 X569-SPLITT-OUT-R-INt 0 X569-SPLITT-OUT-R-IN 0 z0=5 td=9.9ps
X569 X356-LSmitll_SPLITT-OUT-X569-LSmitll_SPLITT-IN X569-LSmitll_SPLITT-OUT-X301-LSmitll_OR2T-INt X569-SPLITT-OUT-R-INt LSmitll_SPLITT

t1810 X570-LSmitll_SPLITT-OUT-X303-LSmitll_OR2T-INt 0 X570-LSmitll_SPLITT-OUT-X303-LSmitll_OR2T-IN 0 z0=5 td=0.7ps
t1811 X570-SPLITT-OUT-R-INt 0 X570-SPLITT-OUT-R-IN 0 z0=5 td=9.8ps
X570 X443-LSmitll_SPLITT-OUT-X570-LSmitll_SPLITT-IN X570-LSmitll_SPLITT-OUT-X303-LSmitll_OR2T-INt X570-SPLITT-OUT-R-INt LSmitll_SPLITT

t1812 X571-LSmitll_SPLITT-OUT-X306-LSmitll_OR2T-INt 0 X571-LSmitll_SPLITT-OUT-X306-LSmitll_OR2T-IN 0 z0=5 td=0.6ps
t1813 X571-SPLITT-OUT-R-INt 0 X571-SPLITT-OUT-R-IN 0 z0=5 td=9.9ps
X571 X343-LSmitll_SPLITT-OUT-X571-LSmitll_SPLITT-IN X571-LSmitll_SPLITT-OUT-X306-LSmitll_OR2T-INt X571-SPLITT-OUT-R-INt LSmitll_SPLITT

t1814 X572-LSmitll_SPLITT-OUT-X310-LSmitll_OR2T-INt 0 X572-LSmitll_SPLITT-OUT-X310-LSmitll_OR2T-IN 0 z0=5 td=0.3ps
t1815 X572-SPLITT-OUT-R-INt 0 X572-SPLITT-OUT-R-IN 0 z0=5 td=10.1ps
X572 X402-LSmitll_SPLITT-OUT-X572-LSmitll_SPLITT-IN X572-LSmitll_SPLITT-OUT-X310-LSmitll_OR2T-INt X572-SPLITT-OUT-R-INt LSmitll_SPLITT

t1816 X573-LSmitll_SPLITT-OUT-X312-LSmitll_OR2T-INt 0 X573-LSmitll_SPLITT-OUT-X312-LSmitll_OR2T-IN 0 z0=5 td=0.8ps
t1817 X573-SPLITT-OUT-R-INt 0 X573-SPLITT-OUT-R-IN 0 z0=5 td=10.3ps
X573 X416-LSmitll_SPLITT-OUT-X573-LSmitll_SPLITT-IN X573-LSmitll_SPLITT-OUT-X312-LSmitll_OR2T-INt X573-SPLITT-OUT-R-INt LSmitll_SPLITT

t1818 X574-LSmitll_SPLITT-OUT-X315-LSmitll_OR2T-INt 0 X574-LSmitll_SPLITT-OUT-X315-LSmitll_OR2T-IN 0 z0=5 td=0.7ps
t1819 X574-SPLITT-OUT-R-INt 0 X574-SPLITT-OUT-R-IN 0 z0=5 td=9.6ps
X574 X351-LSmitll_SPLITT-OUT-X574-LSmitll_SPLITT-IN X574-LSmitll_SPLITT-OUT-X315-LSmitll_OR2T-INt X574-SPLITT-OUT-R-INt LSmitll_SPLITT

t1820 X575-LSmitll_SPLITT-OUT-X320-LSmitll_OR2T-INt 0 X575-LSmitll_SPLITT-OUT-X320-LSmitll_OR2T-IN 0 z0=5 td=1.0ps
t1821 X575-SPLITT-OUT-R-INt 0 X575-SPLITT-OUT-R-IN 0 z0=5 td=10.2ps
X575 X478-LSmitll_SPLITT-OUT-X575-LSmitll_SPLITT-IN X575-LSmitll_SPLITT-OUT-X320-LSmitll_OR2T-INt X575-SPLITT-OUT-R-INt LSmitll_SPLITT

t1822 X576-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-INt 0 X576-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-IN 0 z0=5 td=2.6ps
t1823 X576-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-INt 0 X576-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-IN 0 z0=5 td=3.9ps
X576 GCLK X576-LSmitll_SPLITT-OUT-X423-LSmitll_SPLITT-INt X576-LSmitll_SPLITT-OUT-X524-LSmitll_SPLITT-INt LSmitll_SPLITT

* PTLs from input pads
t876 GCLKt 0 GCLK 0 z0=5 td=17.9ps
t608 program_line4t 0 program_line4 0 z0=5 td=7.0ps
t596 program_line3t 0 program_line3 0 z0=5 td=7.6ps
t588 program_line2t 0 program_line2 0 z0=5 td=5.7ps
t580 program_line1t 0 program_line1 0 z0=5 td=6.0ps
t604 load4t 0 load4 0 z0=5 td=6.0ps
t600 load3t 0 load3 0 z0=5 td=20.7ps
t592 load2t 0 load2 0 z0=5 td=8.4ps
t584 load1t 0 load1 0 z0=5 td=3.1ps

t616 Addr1_1t 0 Addr1_1 0 z0=5 td=11.3ps
t612 Addr1_0t 0 Addr1_0 0 z0=5 td=20.2ps
t624 Addr0_1t 0 Addr0_1 0 z0=5 td=2.6ps
t620 Addr0_0t 0 Addr0_0 0 z0=5 td=14.6ps
t628 read1t 0 read1 0 z0=5 td=6.7ps
t632 read0t 0 read0 0 z0=5 td=11.8ps
t636 read_at_first_addr1t 0 read_at_first_addr1 0 z0=5 td=2.9ps
t640 read_at_first_addr0t 0 read_at_first_addr0 0 z0=5 td=5.5ps

* PTLs to output pads
t1307 bit_out0t 0 bit_out0 0 z0=5 td=18.1ps
t1308 bit_out1t 0 bit_out1 0 z0=5 td=20.0ps
t1309 bit_out2t 0 bit_out2 0 z0=5 td=17.3ps
t1310 bit_out3t 0 bit_out3 0 z0=5 td=19.5ps
t1311 bit_out4t 0 bit_out4 0 z0=5 td=19.6ps
t1312 bit_out5t 0 bit_out5 0 z0=5 td=19.5ps
t1313 bit_out6t 0 bit_out6 0 z0=5 td=17.1ps

.ends programmer_instr_memory_final_route